
//
// TODO: 
//
// 10/10/2018
//
//  - remove loader_checksum as it operates on running_checksum now.
//

//
// See MENLO_COPYRIGHT.TXT for the copyright notice for this file.
//
// Use of this file is not allowed without the copyright notice present
// and re-distributed along with these files.
//

//
// Gigatron BabelFish protocol implemented in System Verilog modeled
// on RDMA.
//
// Normally BabelFish runs on an Arduino, and its source code
// is in the Gigatron Rom Git project at:
//
// https://github.com/kervinck/gigatron-rom/Utils/BabelFish/babelfish.ino
//
// In this case BabelFish is implemented in System Verilog and is
// used by the Gigatron option ROM loader.
//
// Since the BabelFish loader protocol is essentially a version of RDMA
// (Remote Direct Memory Access), it will be modeled as such. This makes
// this Verilog code useful for other projects, such as network connected
// FPGA's for Software Defined Radio (SDR), machine tools (CNC), storage,
// and FPGA assisted high speed network communications between applications.
//
// FUTURE WORK:
//
//  Can generalize this RDMA communications handler by:
//
//  Add an IOMMU module to the output addresses. This will allow
//  address translation, validation, scatter/gather support, as
//  well as translations to program/VM virtual addresses based on
//  platform.
// 
//  Have the link level byte stream module interface be supplied to the
//  RDMA transmitter/receiver rather than contained within. This will allow
//  packet oriented protocols such as ethernet, UDP/IP/TCP to be readily
//  swapped in and out.
//
//  Have the RDMA framer modules interface be provided to the RDMA
//  transmitter/receiver. This allows other formats to be utilized
//  such as Infiniband or system TCP direct data placement.
//

module menlo_babelfish_rdma_transmitter
(
    input fpga_clock,      // FPGA 50Mhz clock
    input gigatron_clock,  // 6.25 Mhz Gigatron clock
    input reset,           // Reset when == 1

    // Timing input from the Gigatron
    input  famicom_pulse, // hsync_n
    input  famicom_latch, // vsync_n

    // Output to the Gigatron generated by this module
    output famicom_data,

    // Signals from user interface to select program to load
    input  request,  // true when user select load
    output request_ack, // true when transfer is complete.

    //
    // This provides access to the program loader option ROM.
    // rom_address == 0 is that start of the GT1 binary program
    // to load, as the invoker handles any translation from the base
    // 0 rom_address here to the offset into the option ROM is required.
    //
    output [15:0] rom_address,
    input [7:0] rom_data
  );

  reg reg_request_ack;
  assign request_ack = reg_request_ack;

  //
  // Current ROM address.
  //
  // This is updated as the state machine walks through the GT1 pages
  // in the option ROM loading them as a series of frames.
  //
  // It provides the base rom address to the frame loader for its
  // data to load. The frame loader will generate its own rom access
  // cycles as required. This register is only updated by this modules state
  // machine.
  //
  reg [15:0] reg_rom_address; // Data address of current program data being loaded.

  // Command to the page loader, and its ack
  reg reg_send_page_request;
  wire send_page_request_ack;

  //
  // The page loaders rom address generation is multiplexed based on
  // whether the page loader is active or not.
  //
  wire [15:0] page_loader_rom_address;

  //
  // This switches the rom address output between this module and
  // the page loader module based on when the page loader is active.
  //
  assign rom_address = (reg_send_page_request == 1'b1) ? page_loader_rom_address : reg_rom_address;

  //
  // The GT1 file loader advances through the ROM starting at address 0
  // reading the series of page headers (address, length), and invoking
  // the page loader for the pages data. The page loader will send the
  // page data as a series of one or more frames and return when done.
  //
  // The last page record in the GT1 file has a high address byte of 0
  // marking the end. The next bytes describe the start address for
  // the program, which is sent as a 0 length page to the page loader,
  // which is an indication to send a single 0 length frame with the
  // start address, as that is the Gigatron loader protocol.
  //

  //
  // At the start of a page send this is the GT1 page address and length.
  //
  // The address here is the remote Gigatron address and length to place
  // the GT1 page to.
  //
  reg [15:0] reg_current_page_remote_address;
  reg [8:0] reg_current_page_remote_length; // must handle 0 - 256 so its 9 bits.

  //
  // Page loader module instance.
  //

  menlo_babelfish_rdma_page_transmitter rdma_page_transmitter (
    .fpga_clock(fpga_clock),
    .gigatron_clock(gigatron_clock),
    .reset(reset),

     // pulse and latch are the input timing control signals.
    .famicom_pulse(famicom_pulse), // input
    .famicom_latch(famicom_latch), // input

    // Data is generated by the loader to be input to the Gigatron
    .famicom_data(famicom_data),  // output

     // These are the page request parameters
    .request(reg_send_page_request),       // input
    .request_ack(send_page_request_ack),   // output

    //
    // This address and length are the values to place in the loader frame
    // to represent the remote page address and length.
    //
    .request_page_remote_address(reg_current_page_remote_address), // input
    .request_page_remote_length(reg_current_page_remote_length),   // input

    //
    // This is the ROM address where the data for the page is.
    // It's length is the reg_current_page_remote_length.
    //
    .request_data_rom_address(reg_rom_address), // input

    // This gives the frame loader access to the option ROM when its active.
    .rom_address(page_loader_rom_address), // output
    .rom_data(rom_data)                   // input
  );

  //
  // GT1 file Loader States:
  //

  parameter[4:0]
    SEND_IDLE             = 5'b00000,

    SEND_FILE             = 5'b00001,

    // Getting Page parameters from the ROM
    PAGE_ADDRESS_HIGH     = 5'b00010,
    PAGE_ADDRESS_LOW      = 5'b00011,
    PAGE_LENGTH           = 5'b00100,

    // Sending a page as a series of frames.
    SENDING_PAGE          = 5'b00101,

    // Send the next page in the ROM.
    SEND_NEXT_PAGE        = 5'b00110,

    // Send a page of the file
    SEND_PAGE             = 5'b00111,

    // Getting the start address page from the ROM
    START_ADDRESS_HIGH    = 5'b01000,

    START_ADDRESS_LOW     = 5'b01001,

    SENDING_START_ADDRESS = 5'b01010,

    SENDING_PAGE_ACK      = 5'b01011,

    // Waiting for the invoker to deassert request and finish.
    FINALIZE              = 5'b11111;

  // Loader state machine
  reg [4:0] loader_state;
  reg [4:0] loader_next_state;

  always@(posedge fpga_clock) begin

    if (reset == 1'b1) begin
      reg_rom_address <= 0;
      reg_request_ack <= 0;

      loader_state <= SEND_IDLE;
      loader_next_state <= SEND_IDLE;

      reg_current_page_remote_address <= 0;
      reg_current_page_remote_length <= 0;

      reg_send_page_request <= 0;
    end
    else begin

      //
      // Not reset
      //

      case (loader_state) 

        SEND_IDLE: begin
          if (request == 1'b1) begin
            reg_request_ack <= 0;
            loader_state <= SEND_FILE;
          end
        end

        SEND_FILE: begin

            //
            // Request to transfer a GT1 file from the start of the ROM
            //
            reg_rom_address <= 0;

            reg_current_page_remote_address <= 0;
            reg_current_page_remote_length <= 0;

            reg_send_page_request <= 0;

            loader_state <= SEND_PAGE;
        end

        SEND_PAGE: begin
            //
            // Current rom_address points to the start byte of the new page
            // which is the high address byte.
            //
            loader_state <= PAGE_ADDRESS_HIGH;
        end

        PAGE_ADDRESS_HIGH: begin

          // Got the remote address high, now get low

          //
          // If its not the first segment of the ROM and the
          // address high byte is 0, then this is the end of
          // the series of segments.
          //
          // The very first segment in the file is allowed to
          // have address high equal to zero in order to support
          // loading varaibles into the zero page.
          // 
          if ((reg_rom_address != 16'h0000) && (rom_data == 8'h00)) begin

            //
            // Address high byte == 0 means end of page records.
            //
            // Next two bytes is the GT1 program start address.
            //
            reg_rom_address <= reg_rom_address + 16'd1;
            loader_state <= START_ADDRESS_HIGH;
          end
          else begin
            // High address byte != 0 and not rom_address == 0, start of new page.
            reg_current_page_remote_address[15:8] <= rom_data;
            reg_rom_address <= reg_rom_address + 16'd1;
            loader_state <= PAGE_ADDRESS_LOW;
          end
        end

        PAGE_ADDRESS_LOW: begin
          // Got the low address, now get the page length
          reg_current_page_remote_address[7:0] <= rom_data;

          // Read the next byte in the ROM
          reg_rom_address <= reg_rom_address + 16'd1;

          loader_state <= PAGE_LENGTH;
        end

        PAGE_LENGTH: begin

          // Got the page length, now send page.

          //
          // Special handling: 0 means 256 bytes in a page.
          //
          // The length is a 9 bit field to accomodate this.
          //
          if (rom_data == 8'h00) begin
            reg_current_page_remote_length <= 9'd256;
          end
          else begin
            reg_current_page_remote_length[8:8] <= 1'b0;
            reg_current_page_remote_length[7:0] <= rom_data;
          end

          // Point to the pages data area in the ROM
          reg_rom_address <= reg_rom_address + 16'd1;

          // Start the page loader, wait for its ack.
          reg_send_page_request <= 1'b1;

          loader_next_state <= SEND_NEXT_PAGE;
          loader_state <= SENDING_PAGE;
        end

        SENDING_PAGE: begin
          // Stay in the SENDING_PAGE state till ack
          if (send_page_request_ack == 1'b1) begin
            reg_send_page_request <= 1'b0;
            loader_state <= SENDING_PAGE_ACK;
          end
        end

        SENDING_PAGE_ACK: begin
          // Wait till ack is deasserted
          if (send_page_request_ack == 1'b0) begin
            loader_state <= loader_next_state;
          end
        end

        SEND_NEXT_PAGE: begin
          // start next page read

          // Advance the  ROM by the data just sent from the current page.
          reg_rom_address <= reg_rom_address + reg_current_page_remote_length;

          loader_state <= SEND_PAGE;
        end

        START_ADDRESS_HIGH: begin
          // High byte of GT1 programs start address.
          reg_current_page_remote_address[15:8] <= rom_data;
          reg_rom_address <= reg_rom_address + 16'd1;
          loader_state <= START_ADDRESS_LOW;
        end

        START_ADDRESS_LOW: begin
          // Low byte of GT1 programs start address
          reg_current_page_remote_address[7:0] <= rom_data;

          //
          // Do not increment the rom address, as we are at the end of the ROM
          // image for this GT1 program.
          //
          //reg_rom_address <= reg_rom_address + 1;

          // Send start address as a parameterized page send of length 0.
          reg_current_page_remote_length <= 9'd0;

          // Start the page loader, wait for its ack.
          reg_send_page_request <= 1'b1;

          loader_next_state <= SENDING_START_ADDRESS;
          loader_state <= SENDING_PAGE;
        end

        SENDING_START_ADDRESS: begin
          // Done with the GT1 file transfer, send ack to invoker.
          reg_request_ack <= 1'b1;

          loader_state <= FINALIZE;
        end

        FINALIZE: begin
          // Stay in finalize state until request is deasserted.
          if (request == 1'b0) begin
            reg_request_ack <= 1'b0;
            loader_state <= SEND_IDLE;
          end
        end

      endcase

    end // not reset

  end // always

  //
  // GT1 File Format:
  //
  // gigatron-rom\Docs\GT1-files.txt
  //
  // The file is sent in frames documented in the babelfish_frame_loader..
  //
  // The file consists of multiple segments with an address,
  // a length, and the bytes. This is because a GT1 program
  // is spread across memory between the video display lines
  // and is how the vCPU executes programs.
  //
  // Each segment can't be any larger than a Gigatron memory
  // page which is 256 bytes. The format represents the maximum
  // length segment as 0, to mean 256 bytes.
  //
  // For the loader, each segment is broken up into one or more transfer
  // frames, each up to 60 bytes.
  //
  // Frames do not cross page (256 byte) boundaries.
  //
  // The end of a series of segments is represented by a high address byte of 0.
  //
  // For this to work, any segment that loads into page 0 must be the first
  // segment in the GT1 file, and only one such segment is allowed. A GT1
  // file with no segments is invalid, so zero handling works.
  //
  // At the end of the series of segments is the program start address
  // as two bytes in high, low order. This is passed in a zero length
  // transfer frame, and an indication its the program start, or go address.
  //
  // see doTransfer() from BabelFish.ino
  //
  // Segment for a specific memory page:
  //
  // Segment X:
  // Byte 0: - address high
  // Byte 1: - address low
  // Byte 2: - length. If 0, its 256.
  // Byte 3: - first data byte
  // Byte x: - last data byte, byte 2 determines length of data.
  // 
  // Segment X + 1:
  // Byte 0: - address high, or 0 if end of segments
  //
  // Last Segment is the GT1 files start address:
  // Byte 0:   - value 0, represents end of series of segments (see above)
  // Byte x:   - start address high
  // Byte x+1: - start address low
  //
  // Note: There is an address overflow check beyond 256 boundary
  // Address Byte 0 if 0 means end of a series of segments. If
  // a pages end address is exceeded, the loader fails.
  //
  // A sendGt1Execute() command is sent to the Gigatron to execute
  // the loaded program. It uses a loader frame with start byte 'L', (0x4C)
  // but a length of 0. The address supplied is the start address.
  //

endmodule // menlo_babelfish_rdma_transmitter

//
// This is the page loader.
//
// It loads the page as a series of frames.
//
// The main BabelFish loader passes the base address of the page
// data in the rom, and the page address and length already read.
//
// Note that a zero length reguest_page_remote_length means
// to send the reguest_page_remote_address as a GT1 program start
// address frame.
//
module menlo_babelfish_rdma_page_transmitter
(
    input fpga_clock,      // FPGA 50Mhz clock
    input gigatron_clock,  // 6.25 Mhz Gigatron clock
    input reset,           // Reset when == 1

    // Timing input from the Gigatron
    input  famicom_pulse,
    input  famicom_latch,

    // Output to the Gigatron generated by this module
    output famicom_data,

    // Signals from invoker
    input  request,     // true when page load is requested
    output request_ack, // true when page load is complete.

    //
    // This address and length are the values to place in the loader frames
    // to represent the remote page address and length.
    //
    input [15:0] request_page_remote_address,
    input [8:0] request_page_remote_length,

    //
    // This is the ROM address where the data for the page is.
    // It's length is the reg_current_page_remote_length.
    //
    input [15:0] request_data_rom_address,

    //
    // This points to the pages data area. Address and length have already
    // been read and passed in as input parameters.
    //
    output [15:0] rom_address,
    input [7:0] rom_data
);

  parameter FRAME_DATA_SIZE = 8'd60;

  reg reg_request_ack;
  assign request_ack = reg_request_ack;

  reg reg_send_frame_request;
  wire send_frame_request_ack;

  //
  // Current ROM address.
  //
  // This is updated as the state machine walks through the data in
  // the page which is sent as a series of frames.
  //
  // It provides the base rom address to the frame loader for its
  // data to load. The frame loader will generate its own rom access
  // cycles as required. This register is only updated by this modules state
  // machine.
  //
  reg [15:0] reg_rom_address; // Data address of current program data being loaded.

  //
  // This is the address output from the frame loader.
  //
  wire [15:0] frame_loader_rom_address;

  //
  // The rom_address is generated by the frame loader. This module
  // does not need to access the rom data directly.
  //
  assign rom_address = frame_loader_rom_address;

  //
  // At the start of a page send this is the GT1 page address and length.
  //
  // The address here is the remote Gigatron address and length to place
  // the GT1 page to.
  //
  // The length is decremented as frames are sent within the page.
  //
  //reg [15:0] reg_current_page_address; // debug
  reg [7:0] reg_current_page_length;

  //
  // This is the address and length that should be sent with the current frame.
  // It does not represent the ROM address, or the GT1 page base address as this
  // must advance with each frames that is a partial GT1 page.
  //
  reg [15:0] reg_current_frame_remote_address;

  // A frame is always 8 bits length, 0 - 60.
  reg [7:0] reg_current_frame_remote_length;

  //
  // This is how much of the current page has been transferred.
  //
  reg [7:0] reg_current_page_length_transferred;

  // total pages sent. Wraps around. For debugging/tracing.
  reg [15:0] reg_total_pages_sent;

  //
  // The running checksum is set at the start of a page
  // and updated by each frame sent.
  //
  // Each frame takes the complement of its current value
  // at the end of the frame and sends that as the frames
  // checksum. If all of the frames bits and previous frames
  // before within the page have been sent ok, then the
  // sum will be zero. Otherwise it indicates a reception
  // error.
  //
  reg [7:0] reg_running_checksum_input;

  //
  // The frame sender provides its updated value of the
  // running checksum at the end of frame send.
  //
  wire [7:0] running_checksum_output;

  //
  // Create an instance of the BabelFish frame loader.
  //
  menlo_babelfish_rdma_frame_transmitter rdma_frame_transmitter (
    .fpga_clock(fpga_clock),
    .gigatron_clock(gigatron_clock),
    .reset(reset),

     // pulse and latch are the input timing control signals.
    .famicom_pulse(famicom_pulse), // input
    .famicom_latch(famicom_latch), // input

    // Data is generated by the loader to be input to the Gigatron
    .famicom_data(famicom_data),  // output

     // These are the frame request parameters
    .request(reg_send_frame_request),       // input
    .request_ack(send_frame_request_ack),   // output

    //
    // This address and length are the values to place in the loader frame
    // to represent the remote page address and length.
    //
    .request_frame_remote_address(reg_current_frame_remote_address), // input
    .request_frame_remote_length(reg_current_frame_remote_length),   // input

    //
    // This is the ROM address where the data for the frame is.
    // It's length is the request_frame_remote_length.
    //
    .request_data_rom_address(reg_rom_address), // input

    // This gives the frame loader access to the option ROM when active.
    .rom_address(frame_loader_rom_address), // output
    .rom_data(rom_data),        // input

    //
    // Frame sender receives the running checksum at start,
    // and outputs its new value at end.
    //
    .running_checksum_input(reg_running_checksum_input),
    .running_checksum_output(running_checksum_output)

  );

  //
  // BabelFish GT1 page loader state machine.
  //

  //
  // Loader States:
  //

  parameter[3:0]
    SEND_IDLE             = 4'b0000,

    // Send a page of the file
    SEND_PAGE             = 4'b0001,

    // Send a page consisting as one or more frames
    SENDING_PAGE_FRAMES   = 4'b0010,

    // Send page is complete
    SEND_PAGE_COMPLETE    = 4'b0011,

    SEND_START_ADDRESS    = 4'b0100,

    SENDING_START_ADDRESS = 4'b0101,

    // Sending a frame within a page
    SENDING_FRAME         = 4'b0110,

    // Frame send completed
    SENDING_FRAME_ACK     = 4'b0111,

    // Waiting for the invoker to deassert request and finish.
    FINALIZE              = 4'b1000;

  // Loader state machine
  reg [3:0] loader_state;
  reg [3:0] loader_next_state;

  always@(posedge fpga_clock) begin

    if (reset == 1'b1) begin
      reg_rom_address <= 0;
      reg_request_ack <= 0;
      reg_send_frame_request <= 0;

      loader_state <= SEND_IDLE;
      loader_next_state <= SEND_IDLE;

      reg_total_pages_sent <= 0;

      //reg_current_page_address <= 0;
      reg_current_page_length <= 0;
      reg_current_frame_remote_address <= 0;
      reg_current_frame_remote_length <= 0;
      reg_current_page_length_transferred <= 0;

      reg_running_checksum_input <= 0;
    end
    else begin

      //
      // Not reset
      //

      case (loader_state) 

        SEND_IDLE: begin
          if (request == 1'b1) begin

            reg_request_ack <= 0;

            //
            // Request to transfer a GT1 page from the ROM.
            //

            //
            // Load control variables from the parameters.
            //
            //reg_current_page_address <= request_page_remote_address;

            reg_current_page_length <= request_page_remote_length[7:0];

            // First frame of the page.
            reg_current_frame_remote_address <= request_page_remote_address;

            reg_rom_address <= request_data_rom_address;
            reg_current_frame_remote_address <= request_page_remote_address;

            // This is only 8 bits for each frame is 0 - 60.
            reg_current_frame_remote_length <= request_page_remote_length[7:0];

            reg_current_page_length_transferred <= 0;

            reg_total_pages_sent <= reg_total_pages_sent + 16'd1;

            //
            // Initialize the running checksum to 'g' (0x67)
            //
            reg_running_checksum_input <= 8'h67;

            if (request_page_remote_length == 9'd0) begin
              // Request to send start address frame.
              loader_state <= SEND_START_ADDRESS;
            end
            else begin
              // Send a data page.
              loader_state <= SEND_PAGE;
            end
          end
        end

        SEND_PAGE: begin

          if (reg_current_page_length > FRAME_DATA_SIZE) begin
              // Must send page in multiple frames
              reg_current_frame_remote_length <= FRAME_DATA_SIZE;

              // Set the amount transferred to the size of the first frame
              reg_current_page_length_transferred <= FRAME_DATA_SIZE;

              // Decrement the bytes left in the page.
              reg_current_page_length <= reg_current_page_length - FRAME_DATA_SIZE;
          end
          else begin
              reg_current_frame_remote_length <= reg_current_page_length;

              // Set the amount transferred to the size of the first frame
              reg_current_page_length_transferred <= reg_current_page_length;

              // Last frame in the page.
              reg_current_page_length <= 0;
          end

          // Send frame
          reg_send_frame_request <= 1'b1;

          loader_next_state <= SENDING_PAGE_FRAMES;
          loader_state <= SENDING_FRAME;
        end

        SENDING_PAGE_FRAMES: begin

          //
          // Update the current rom address and the page remote address with
          // what was just transferred in the last frame.
          //
          reg_rom_address <= reg_rom_address + reg_current_frame_remote_length;

          reg_current_frame_remote_address <= reg_current_frame_remote_address + 
                                              reg_current_frame_remote_length;

          //
          // Update the running checksum with the value from the frame.
          //
          reg_running_checksum_input <= running_checksum_output;

          if (reg_current_page_length == 8'h00) begin
            // Done
            loader_state <= SEND_PAGE_COMPLETE;
          end
          else begin
            // Send next frame in the page
            if (reg_current_page_length > FRAME_DATA_SIZE) begin
              reg_current_frame_remote_length <= FRAME_DATA_SIZE;

              // Update total transferred
              reg_current_page_length_transferred <= reg_current_page_length_transferred + FRAME_DATA_SIZE;

              reg_current_page_length <= reg_current_page_length - FRAME_DATA_SIZE;
            end
            else begin
              reg_current_frame_remote_length <= reg_current_page_length;

              reg_current_page_length_transferred <= reg_current_page_length_transferred +
                                                     reg_current_page_length;

              // Last frame
              reg_current_page_length <= 0;
            end

            // Send next frame
            reg_send_frame_request <= 1'b1;

            loader_next_state <= SENDING_PAGE_FRAMES;
            loader_state <= SENDING_FRAME;
          end // not done loading page
        end

        SEND_PAGE_COMPLETE: begin
          // Ackknowledge we are done
          reg_request_ack <= 1'b1;

          loader_state <= FINALIZE;
        end

        SEND_START_ADDRESS: begin

          // Send 0 length frame
          reg_send_frame_request <= 1'b1;

          loader_next_state <= SENDING_START_ADDRESS;
          loader_state <= SENDING_FRAME;
        end

        SENDING_START_ADDRESS: begin

          //
          // sending start address frame that defines the GT1 programs entry.
          //

          // Done, ack the invoker
          reg_request_ack <= 1'b1;
          loader_state <= FINALIZE;
        end

        SENDING_FRAME: begin
          // Stay in the SENDING_FRAME state till ack
          if (send_frame_request_ack == 1'b1) begin
            reg_send_frame_request <= 1'b0;
            loader_state <= SENDING_FRAME_ACK;
          end
        end

        SENDING_FRAME_ACK: begin
          // Wait till ack is deasserted
          if (send_frame_request_ack == 1'b0) begin
            loader_state <= loader_next_state;
          end
        end

        FINALIZE: begin
          // Stay in finalize state until request is deasserted.
          if (request == 1'b0) begin
            reg_request_ack <= 1'b0;
            loader_state <= SEND_IDLE;
          end
        end

        default: begin
          loader_state <= SEND_IDLE;
        end

      endcase

    end // not reset

  end // always

endmodule // menlo_babelfish_rdma_page_transmitter

//
// Gigatron RDMA frame transmitter.
//
// A Gigatron loader frame consits of up to 518 bits sent during a
// VSYNC interval, clocked by HSYNC.
//
// The frame contains the remote Gigatron load address, a 6 bit length, and up to
// 60 bytes of data and a checksum.
//
// A frame length of 0 indicates that a start program address frame should
// be sent.
//
module menlo_babelfish_rdma_frame_transmitter
(
    input fpga_clock,      // FPGA 50Mhz clock
    input gigatron_clock,  // 6.25 Mhz Gigatron clock
    input reset,           // Reset when == 1

    // pulse and latch are the input timing control signals.
    input  famicom_pulse,  // hsync_n
    input  famicom_latch,  // vsync_n

    // Data is generated by the loader to be input to the Gigatron
    output famicom_data,

    // Parameters from main BabelFish loader state machine.
    input  request,     // frame send request
    output request_ack, // frame send done.

    //
    // This address and length are the values to place in the loader frame
    // to represent the remote page address and length.
    //
    input [15:0] request_frame_remote_address,
    input [7:0] request_frame_remote_length,

    //
    // This is the ROM address where the data for the frame is.
    // It's length is the request_frame_remote_length.
    //
    input [15:0] request_data_rom_address,

    // These are the signals to read bytes from the ROM
    output [15:0] rom_address,
    input [7:0] rom_data,

    //
    // running_checksum_input is the current running
    // checksum at the start of the frame.
    //
    input [7:0]  running_checksum_input,

    //
    // running_checksum_output is the final calculated
    // checksum when the frame send has completed.
    //
    output [7:0] running_checksum_output
);

  reg reg_request_ack;
  assign request_ack = reg_request_ack;

  reg [15:0] reg_rom_address; // Data address of current program data being loaded.
  assign rom_address = reg_rom_address;

  reg [7:0] reg_running_checksum_output;
  assign running_checksum_output = reg_running_checksum_output;

  // Running checksum of the current frame
  reg [7:0] loader_checksum;

  // Set when in loader mode
  //reg       reg_loader_active; // debug

  //
  // This indicates when bits are to be sent, the parameters, and the ack.
  //
  reg reg_send_bits_request;
  reg reg_send_bits_frame_start;
  reg [7:0] reg_send_bits_value;
  reg [3:0] reg_send_bits_count;

  wire send_bits_request_ack;

  //
  // Loader States:
  //
  // Unlike C code in which the sequence is contained in the order
  // of the source lines, Verilog/FPGA's must explicitly encode
  // the states. This is very similar to async programming in device
  // drivers, but in this case its every single clock cycle.
  //

  // rdma_frame_transmitter states
  parameter[3:0]
    SEND_IDLE             = 4'b0000,
    SENDING_START         = 4'b0001, // (command byte) // 8 bits 'L' (0x4C)
    SENDING_LENGTH        = 4'b0010, // 6 bits
    SENDING_ADDRESS_HIGH  = 4'b0011, // 8 bits
    SENDING_ADDRESS_LOW   = 4'b0100, // 8 bits
    SENDING_DATA          = 4'b0101, // rom_length 8 bit data bytes
    SENDING_CHECKSUM      = 4'b0110, // 8 bits
    SENDING_BYTE          = 4'b0111,
    WAITING_FOR_ACK_N     = 4'b1000,
    SEND_BYTE_FROM_ROM    = 4'b1001,
    READING_BYTE_FROM_ROM = 4'b1010,
    BYTE_READ_FROM_ROM    = 4'b1011,
    FINALIZE              = 4'b1100,
    ADDING_START_CHECKSUM = 4'b1101,
    ADDING_START_CHECKSUM2 = 4'b1110;

  // Loader state machine
  reg [3:0] loader_state;
  reg [3:0] loader_next_state;

  reg [7:0] reg_data_to_transfer;

  // total frames sent. Wraps around. For debugging/tracing.
  reg [15:0] reg_total_frames_sent;

  //
  // Bit sender subsystem.
  //
  menlo_babelfish_rdma_linklayer_byte_transmitter rdma_byte_transmitter (
    .fpga_clock(fpga_clock),
    .reset(reset),
    .value(reg_send_bits_value),
    .number_of_bits(reg_send_bits_count),
    .pulse(famicom_pulse),          // hsync_n, famicom_pulse
    .latch(famicom_latch),          // vsync_n, famicom_latch
    .frame_start(reg_send_bits_frame_start),    // set if this is the first byte of the frame.
    .output_port(famicom_data),     // famicom_data
    .request(reg_send_bits_request),
    .request_ack(send_bits_request_ack)
  );

  // Debug
  //reg debug_transmitting_checksum; // debug

  always@(posedge fpga_clock) begin

    if (reset == 1'b1) begin
      reg_request_ack <= 0;
      //reg_loader_active <= 0;

      loader_state <= SEND_IDLE;
      loader_next_state <= SEND_IDLE;

      loader_checksum <= 0;

      reg_running_checksum_output <= 0;

      reg_rom_address <= 16'h0;
      reg_data_to_transfer <= 0;

      reg_total_frames_sent <= 0;

      //
      // communication variable with the send bits process.
      //
      reg_send_bits_request <= 1'b0;
      reg_send_bits_frame_start <= 1'b0;
      reg_send_bits_value <= 8'b0;
      reg_send_bits_count <= 4'b0;

      // Debug
      //debug_transmitting_checksum <= 0;

    end
    else begin

      //
      // Not reset
      //

      case (loader_state) 

        SEND_IDLE: begin

          if (request == 1'b1) begin

            //debug_transmitting_checksum <= 1'b0;

            //
            // Transfer the current running checksum input
            // to the local running checksum register.
            //
            reg_running_checksum_output <= running_checksum_input;

            //
            // Request to transfer a frame.
            //
            reg_request_ack <= 0;
            //reg_loader_active <= 1'b1;

            // Send first byte with frame_start attribute
            reg_send_bits_value <= 8'h4C; // start byte 'L'

            // Set rom address to 0 which points to start of the data.
            reg_rom_address <= 16'h0;

            reg_send_bits_count <= 4'd8;

            //
            // This is the start of a frame. This has the byte
            // transmitter wait a vsync_n cycle from LOW => HIGH => LOW.
            //
            reg_send_bits_frame_start <= 1'b1;

            reg_total_frames_sent <= reg_total_frames_sent + 16'd1;

            //
            // Note: Addition to the checksum for the frame start
            // handling must occur over multiple clock cycles
            // since the Verilog statements only allow one assignment
            // and result per clock cycle. A parallel implementation
            // could be used, but we have time here do to this
            // before the next vsync_n cycle.
            //
            // Yes, we are starting with constants here, but the
            // receiver will not, so the code is similar. Plus this
            // module could be used in the future with different
            // start bytes as a parameter to support Gigatron keyboard
            // and command input.
            //

            //
            // Checksum starts with 'g' 0x67.
            //
            loader_checksum <= 8'h67;

            // Must frame start byte to checksum before send.
            loader_state <= ADDING_START_CHECKSUM;
          end
        end

        ADDING_START_CHECKSUM: begin

          //
          // Current byte being sent is pre-added to the running
          // checksum.
          //

          loader_checksum <= loader_checksum + 8'h4C;

          reg_running_checksum_output <= reg_running_checksum_output + 8'h4C;

          loader_state <= ADDING_START_CHECKSUM2;
        end

        ADDING_START_CHECKSUM2: begin

          //
          // Note: Gigatron's BabelFish.ino also shifts the frame
          // start byte left by 6 and adds it to the checksum again.
          //
          loader_checksum <= loader_checksum + (8'h4C << 6);

          reg_running_checksum_output <= reg_running_checksum_output + 
            (8'h4C << 6);

          // Start the byte transmission sequence
          reg_send_bits_request <= 1'b1;

          // return to SENDING_START state when done
          loader_next_state <= SENDING_START;

          // In SENDING_BYTE state
          loader_state <= SENDING_BYTE;

        end

        SENDING_START: begin

          //
          // sending start byte has completed, this is not set for
          // the rest of the bytes.
          //
          reg_send_bits_frame_start <= 1'b0;

          // Send frame data length byte passed from the invoker
          reg_send_bits_value <= request_frame_remote_length;

          // Length is sent as 6 bits in the frame protocol.
          reg_send_bits_count <= 4'd6;

          loader_checksum <= loader_checksum + request_frame_remote_length;

          reg_running_checksum_output <= reg_running_checksum_output + 
            request_frame_remote_length;

          reg_send_bits_request <= 1'b1;

          loader_next_state <= SENDING_LENGTH;
          loader_state <= SENDING_BYTE;
        end

        SENDING_LENGTH: begin

          //
          // sending length byte has completed
          //

          // The rest of the byte transfers in the frame will be 8 bit.
          reg_send_bits_count <= 4'd8;

          // Send the high address byte
          reg_send_bits_value <= request_frame_remote_address[15:8];

          // Keep checksum updated with current byte being sent.
          loader_checksum <= loader_checksum + request_frame_remote_address[15:8];

          reg_running_checksum_output <= reg_running_checksum_output +
            request_frame_remote_address[15:8];

          reg_send_bits_request <= 1'b1;

          loader_next_state <= SENDING_ADDRESS_HIGH;
          loader_state <= SENDING_BYTE;
        end

        SENDING_ADDRESS_HIGH: begin

          // Send the low address byte
          reg_send_bits_value <= request_frame_remote_address[7:0];

          // Keep checksum updated with current byte being sent.
          loader_checksum <= loader_checksum + request_frame_remote_address[7:0];

          reg_running_checksum_output <= reg_running_checksum_output +
            request_frame_remote_address[7:0];

          reg_send_bits_request <= 1'b1;

          loader_next_state <= SENDING_ADDRESS_LOW;
          loader_state <= SENDING_BYTE;
        end

        SENDING_ADDRESS_LOW: begin

          // Set data start address to the ROM
          reg_rom_address <= request_data_rom_address;

          //
          // request_frame_remote_length is the total data length
          // to transfer.
          //
          // It uses 0 to indicate the sending of a program address start frame.
          // In this case no data payload is sent, just the ending checksum.
          //
          if (request_frame_remote_length == 8'h00) begin

              // There are no data bytes to send. Send the checksum and complete.
              reg_data_to_transfer <= 8'h00;

              loader_state <= SENDING_DATA;
          end
          else begin

              //
              // Set the data to be transferred count, subtract one to
              // account for the first byte sent.
              //
              reg_data_to_transfer <= request_frame_remote_length - 8'd1;

              //
              // Transfer the byte from the ROM.
              //
              // The SEND_BYTE_FROM_ROM state machine keeps the running
              // loader_checksum updated with each data bytes sent.
              //
              loader_next_state <= SENDING_DATA;
              loader_state <= SEND_BYTE_FROM_ROM;
          end
        end

        SENDING_DATA: begin

          if (reg_data_to_transfer == 8'h00) begin

              // Done with data transfer, send the checksum
              //debug_transmitting_checksum <= 1'b1;

              // TODO: validating
              //reg_send_bits_value <= loader_checksum;

              //
              // This math has been validated to be the
              // two's complement of the running checksum.
              //
              // The running checksums complement is sent.
              reg_send_bits_value <= 8'd0 - reg_running_checksum_output;

              reg_send_bits_request <= 1'b1;

              loader_next_state <= SENDING_CHECKSUM;
              loader_state <= SENDING_BYTE;
          end
          else begin

              //
              // Transfer the next data byte from the ROM.
              // It updates the checksum with the data bytes value.
              //

              // Advance the ROM address to the next byte to send.
              reg_rom_address <= rom_address + 16'd1;

              // Decrement the transfer count for this byte being sent.
              reg_data_to_transfer <= reg_data_to_transfer - 8'd1;

              // Stay in SENDING_DATA state until all data bytes sent
              loader_next_state <= SENDING_DATA;
              loader_state <= SEND_BYTE_FROM_ROM;
          end
        end

        SENDING_CHECKSUM: begin

          //
          // Done with frame, send ack to invoker.
          //
          reg_request_ack <= 1'b1;

          //reg_loader_active <= 1'b0;

          // Finalize waits for request to deassert
          loader_state <= FINALIZE;
        end

        FINALIZE: begin

          // Stay in finalize state until request is deasserted.
          if (request == 1'b0) begin
            reg_request_ack <= 1'b0;
            loader_state <= SEND_IDLE;
          end

        end

        //
        // Reading a byte from the ROM and then sending it to the
        // babelfish_bit_sender is a common operation used for
        // each byte in the frame envelope, so make it a common
        // state machine.
        //

        SEND_BYTE_FROM_ROM: begin

          //
          // reg_rom_address has been set
          //
          // loader_next_state has been set by invoker.
          //
          // This entry gives 1 clock to access ROM from when the
          // rom_address was set by the invoker.
          //
          loader_state <= READING_BYTE_FROM_ROM;
        end

        READING_BYTE_FROM_ROM: begin

          // byte to send is in the rom_data.
          reg_send_bits_value <= rom_data;

          // reg_send_bits_count is set by the invoker

          // Update the checksum with the data byte from the ROM
          loader_checksum <= loader_checksum + rom_data;

          reg_running_checksum_output <= reg_running_checksum_output + rom_data;

          // next clock will have data in send_bits_value register
          loader_state <= BYTE_READ_FROM_ROM;
        end

        BYTE_READ_FROM_ROM: begin
          // Now send the byte to the bit sender
          reg_send_bits_request <= 1'b1;
          loader_state <= SENDING_BYTE;
        end

        //
        // Each byte sent uses the following two states to handle
        // hand shake with the babelfish_bit_sender module.
        //
        // loader_next_state is used to return to the previous transfer
        // phase when done.
        //

        SENDING_BYTE: begin
          // Sending byte. Wait for ACK
          if (send_bits_request_ack == 1'b1) begin
            // Request has acknowledged, deassert request, wait for ack to drop.
            reg_send_bits_request <= 1'b0;
            loader_state <= WAITING_FOR_ACK_N;
          end
        end

        WAITING_FOR_ACK_N: begin
          if (send_bits_request_ack == 1'b0) begin
            // ack has dropped.

            // loader_next_state was set by state sending the byte.
            loader_state <= loader_next_state;
          end
        end

        default: begin
          loader_state <= SEND_IDLE;
        end

      endcase

    end

  end // always

  //
  // The Gigatron/BabelFish frame protocol is as follows:
  //
  // A bit stream of 518 total bits.
  //
  // Start of the bitstream is clocked by gigatron_famicom_latch (vsync_n) going high.
  //
  // Each bit is clocked by gigatron_famicom_pulse (hsync_n) going high.
  //
  // The bit is placed on gigatron_famicom_data as input to the Gigatron.
  // 
  // Order sent:
  //
  // Note: all bits are sent MSB first.
  //
  // 8 bits - start byte 'L' (0x4C)
  // 6 bits - block_length
  // 8 bits - address_high
  // 8 bits - address_low
  // 8 bits - data_byte[0]
  // 8 bits - data_byte [block_length - 1]
  // 8 bits - checksum
  //
  
  //
  // Note: There is a place where (2) bits are dropped on purpose
  // due to Gigatron loader timings. Ensure this is implemented
  // in the state machine above. It shows up in the (6) bit
  // length period.
  //

endmodule // menlo_babelfish_rdma_frame_transmitter

//
// Gigatron RDMA byte transmitter.
//
// latch is the vsync_n signal from the Gigatron which indicates
// the start of the frame to send.
//
// pulse is the hsync_n signal from the Gigatron which times
// the bit send rate.
//
// frame_start is set for the first byte of the frame and syncs
// with vsync_n (latch) and hsync_h (pulse) for the sending of
// the first byte before sending the rest of the frame. It should
// only be set for the first byte of the frame, and only the first
// bit will perfom the protocols specific synchronization.
//
// Bits are sent MSB first, up to number_of_bits.
//
// Request handshake protocol:
//
// Note that this is used by each module.
//
// Invoker: (The module requesting service from this module)
//
// Reset starts with request, and request_ack == 1'b0.
//
// Invoker sets request == 1'b1, and waits until request_ack
// becomes 1'b1.
//
// Invoker de-asserts request by setting it to 1'b0, and waits
// until request_ack becomes == 1'b0 before asserting a new request
// again for at least a one clock delay to ensure the de-assertion
// is observed by receiver.
//
// Receiver: (the module implementing the receiver)
//
// Receiver starts with request and request_ack == 1'b0 and
// internally in the IDLE state.
//
// Receiver when in IDLE state receives request == 1'b1, and sets
// an internal register to latch the request. It then performs the
// request asynchronously based on its internal state machine.
//
// When the request is complete it sets request_ack == 1'b1, and
// then goes into a state to await the de-assertion of request to 1'b0.
//
// When request becomes 1'b0, it clears request_ack and goes back
// to the idle state to begin await a new request.
//
module menlo_babelfish_rdma_linklayer_byte_transmitter (
  input fpga_clock,
  input reset, // high true
  input [7:0] value,
  input [3:0] number_of_bits,
  input pulse,          // hsync_n, famicom_pulse
  input latch,          // vsync_n, famicom_latch
  input frame_start,    // set if this is the first byte of the frame.
  output output_port,   // famicom_data
  input  request,
  output request_ack
  );

  reg reg_output_port;
  assign output_port = reg_output_port;

  reg reg_request_ack;
  assign request_ack = reg_request_ack;

  reg [7:0] reg_send_bits_value;

  // total bytes sent. Wraps around. For debugging/tracing.
  reg [15:0] reg_total_bytes_sent;

  // rdma_byte_transmitter states
  parameter[2:0]
    BITS_IDLE               = 3'b000,
    BITS_TRANSFER_NEXT_BIT  = 3'b001,
    BITS_WAIT_H_PULSE_LOW   = 3'b010,
    BITS_WAIT_H_PULSE_HIGH  = 3'b011,
    BITS_WAIT_V_LATCH_LOW   = 3'b100,
    BITS_WAIT_V_LATCH_HIGH  = 3'b101,
    BITS_SENDING_ACK        = 3'b110,
    BITS_UNASSIGNED         = 3'b111;

  reg [2:0] bits_state;

  // Bits are sent MSB first, so this counts down.
  reg [3:0] reg_bits_counter;

  always@(posedge fpga_clock) begin

    if (reset == 1'b1) begin
      bits_state <= BITS_IDLE;
      reg_request_ack <= 1'b0;
      reg_send_bits_value <= 0;
      reg_bits_counter <= 0;

      reg_total_bytes_sent <= 0;

      // This is the data out to the Gigatron's input port bit
      reg_output_port <= 0;
    end
    else begin

      //
      // Not reset
      //

      case (bits_state) 

        BITS_IDLE: begin

          if (request == 1'b1) begin

            //
            // Command to send bits in value, count registers.
            //
            reg_send_bits_value <= value;

            reg_total_bytes_sent <= reg_total_bytes_sent + 16'd1;

            //
            // Send starts at bit 7 (MSB) for 8 bits
            // and bit 5 (MSB) for 6 bits transfer.
            //
            reg_bits_counter <= number_of_bits - 4'd1;

            if (frame_start == 1'b1) begin

              //
              // Protocol:
              //
              // First bit of first byte syncs with VSYNC for start of frame.
              //
              // Frame start sequence:
              //
              // 1) wait for vsync_n to be HIGH
              //
              // 2) Drive first bit onto output port
              //
              // 3) wait for vsync_n going LOW (negative edge)
              //
              // Note: At his point its the normal per bit handshake
              // with hsync_n.
              //
              // 4) wait for hsync_n to be LOW
              //
              // 5) wait for hsync_n to be HIGH (positive edge)
              //
              // 6) send rest of 7 bits using normal per bit handshake.
              //

              bits_state <= BITS_WAIT_V_LATCH_HIGH;
            end
            else begin
              bits_state <= BITS_TRANSFER_NEXT_BIT;
            end
          end
        end

        BITS_TRANSFER_NEXT_BIT: begin

          //
          // Protocol:
          //
          // Transfer a bit.
          //
          // bits are transfered with the following sequence:
          //
          // A) bit is set on the output port
          //
          // B) wait for hsync_n to be LOW
          //
          // C) wait for hsync_n to be HIGH (posedge)
          //     - receiver samples the bit at the HIGH positive edge.
          //

          //
          // Bit send state #A
          //
          // reg_bits_counter contains the index of the current
          // bit to send from 7 - 0. It counts down as the protocol
          // sends MSB first.
          //
          // Note end is underflow wrap around since bit 0 in the count down
          // must be sent before terminating.
          //
          if (reg_bits_counter != 4'b1111) begin
            reg_output_port <= reg_send_bits_value[reg_bits_counter];
            bits_state <= BITS_WAIT_H_PULSE_LOW;
          end
          else begin
            reg_request_ack <= 1'b1;
            bits_state <= BITS_SENDING_ACK;
          end
        end

        BITS_WAIT_H_PULSE_LOW: begin

          //
          // Bit send state #B
          //
          // Waiting for hsync_n to be LOW
          //
          if (pulse == 1'b0) begin
            bits_state <= BITS_WAIT_H_PULSE_HIGH;
          end
        end

        BITS_WAIT_H_PULSE_HIGH: begin

          //
          // Bit send state #C
          //
          // Waiting for hsync_n to be HIGH
          //
          if (pulse == 1'b1) begin

            // Current bit transfer has completed, update the counter.
            reg_bits_counter <= reg_bits_counter - 4'd1;

            bits_state <= BITS_TRANSFER_NEXT_BIT;
          end
        end

        BITS_WAIT_V_LATCH_HIGH: begin

          //
          // In frame start sequence state #1
          //
          // Waiting for vsync_n latch signal to be high which
          // starts the frames sequence.
          //
          if (latch == 1'b1) begin

            //
            // vsync_n is high, transfer first bit and wait for vsync_n == low
            //
            // Frame start sequence state #2
            //
            reg_output_port <= reg_send_bits_value[reg_bits_counter];

            bits_state <= BITS_WAIT_V_LATCH_LOW;
          end
        end

        BITS_WAIT_V_LATCH_LOW: begin

          //
          // In frame start sequence state #3
          //
          // Waiting for vsync_n latch signal to be low
          //
          if (latch == 1'b0) begin

            //
            // To complete the start sequence:
            //
            // 4) wait for hsync_n to be LOW
            //
            // 5) wait for hsync_n to be HIGH
            //
            // 6) send rest of 7 bits using normal per bit handshake.
            //

            //
            // Finish the hsync_n synchronization and then transfer the
            // rest of the 7 bits normally.
            //

            // Transfer the rest of the bits normally on each pulse from hsync_n.
            bits_state <= BITS_WAIT_H_PULSE_LOW;
          end
        end

        BITS_SENDING_ACK: begin

          //
          // Waiting for request to be de-asserted
          //
          if (request == 1'b0) begin
            reg_request_ack <= 1'b0;
            bits_state <= BITS_IDLE;
          end

        end

        default: begin
          bits_state <= BITS_IDLE;
        end

      endcase

    end // not reset

  end // always sendBits

  // 
  // Protocol:
  //
  // From https://github.com/kervinck/gigatron-rom/Utils/BabelFish/babelfish.ino
  //
  // void sendFirstByte(byte value)
  // {
  //   //
  //   // Wait vertical sync NEGATIVE edge to sync with loader
  //   //
  //
  //   // Ensure vSync is HIGH first
  //   while (~PINB & gigatronLatchBit)
  //     ;
  // 
  //   // Send first bit in advance
  //   if (value & 128)
  //     PORTB |= gigatronDataBit;
  //   else
  //     PORTB &= ~gigatronDataBit;
  // 
  //   // Then wait for vSync to drop
  //   while (PINB & gigatronLatchBit)
  //     ;
  // 
  //   //
  //   // Wait for bit transfer at horizontal sync RISING edge. As this is at
  //   // the end of a short (3.8 us) pulse following VERY shortly (0.64us) after
  //   // vSync drop, this timing is tight. That is the reason that interrupts
  //   // must be disabled on the microcontroller and that 1 MHz is not enough.
  //   //
  //   while (PINB & gigatronPulseBit) // Ensure hSync is LOW first
  //     ;
  //   while (~PINB & gigatronPulseBit) // Then wait for hSync to rise
  //     ;
  // 
  //   // Send remaining bits
  //   sendBits(value, 7);
  // }
  // 
  // Send n bits, highest first
  // void sendBits(byte value, byte n)
  // {
  //   for (byte bit=1<<(n-1); bit; bit>>=1) {
  //     // Send next bit
  //     if (value & bit)
  //       PORTB |= gigatronDataBit;
  //     else
  //       PORTB &= ~gigatronDataBit;
  // 
  //
  //     //
  //     // Wait for bit transfer at horizontal sync POSITIVE edge.
  //     //
  //
  //     // Ensure hSync is LOW first
  //     while (PINB & gigatronPulseBit)
  //       ;
  //
  //     // Then wait for hSync to rise
  //     while (~PINB & gigatronPulseBit)
  //       ;
  //   }
  //
  //   // Note: This is handled by the invoker for the Verilog implementation here.
  //   checksum += value;
  // }
  // 
  // Send execute command
  //
  // void sendGt1Execute(word address, byte data[])
  // {
  //   critical();
  //   resetChecksum();
  //   sendFrame('L', 0, address, data);
  //   nonCritical();
  // }
  //

endmodule // menlo_babelfish_rdma_byte_transmitter

//
// Gigatron RDMA Receiver.
//
// The Gigatron loader protocol is a form of RDMA, otherwise known
// as Remote Direct Memory Access. As such, this will be modeled as
// a specific variation/implementation of the general RDMA protocol
// pattern. This will make this logic useful in other projects, such
// as RDMA over ethernet/UDP/IP for SDR radios (Software Defined Radio).
//
// As an RDMA protocol, the receiver just sees a series of receive data
// frames with the address, length, and data to deposit into memory.
//
// The memory is addressed through the passed in RAM signals, allowing
// direct addressing of the RAM. The address range of this RAM must
// accommodate the address ranges of the received RDMA frames.
//
// Currently no out of range checking is done, but a caller
// could limit the memory view port visibility to contain
// a transfer, or remap it similar to an IOMMU handling a scatter/gather
// list and validating for out of range memory accesses.
//
// Such inward DMA mapping and validation would be based on caller
// managed client context, or flow, which would DMA only to
// pre-authorized memory locations.
//
// This support is out of scope for this level, and would be
// provided by a higher level memory and transfer management module.
//
// Details on the Gigatron BabelFish Implementation:
//
// Receive a set of memory pages from a remote system over
// a serial bit stream clocked by the vsync_n and hsync_n
// sync pulses.
//
// The per page data is sent as a series of serial frames containing
// the address, length, and data to be deposited into memory from
// the frame. This is accomplished through the ram_address, ram_data,
// ram_write signals.
//
// At the end, a 0 length frame is received which contains the
// program start address, which is returned separately.
//
// Unlike the menlo_babelfish_transmitter, there is no page handler
// in the receiver chain because the pages are a loader file/ROM format
// unseen by the receiver and all that are scene here are RDMA frames.
//
// The transmission is terminated by the receipt of the start address frame.
//
// The start address received is returned.
//
// Reception commences when the first frame with a valid checksum
// is received after a vsync_n pulse going high. Reception of frames
// continues at each vsync_n going high until the recept of the start
// address frame, or an error from the lower protocol.
//
// If error, this error is returned.
//
// On success, the received start address is returned so that
// the program may be executed.
//
module menlo_babelfish_rdma_receiver (

    input fpga_clock,      // FPGA 50Mhz clock
    input gigatron_clock,  // 6.25 Mhz Gigatron clock
    input reset,           // Reset when == 1

    // pulse and latch are the input timing control signals.
    input  famicom_pulse, // hsync_n
    input  famicom_latch, // vsync_n

    // Serial data input
    input  famicom_data,

    // request/ack signals
    input  request,
    output request_ack,

    // This is the received program start address.
    output [15:0] start_address,

    //
    // This is a real time indication of the receiver state.
    //
    // bits [3:0] frame state.
    // bits [7:5] bit serializer state.
    //
    output [7:0]  receiver_realtime_state,

    // Receive error, and diagnostic state
    output        receive_error,
    output [7:0]  receive_error_state,

    output [15:0] ram_address,
    output [7:0]  ram_data,
    output        ram_write
  );

  reg reg_request_ack;
  assign request_ack = reg_request_ack;

  reg reg_receive_error;
  assign receive_error = reg_receive_error;

  reg [4:0] reg_receive_error_state;
  assign receive_error_state[4:0] = reg_receive_error_state;
  assign receive_error_state[7:5] = 3'b000;

  // This is the output from the frame receiver
  wire [4:0] frame_receiver_error_state;

  reg reg_receive_frames_request;
  wire receive_frames_request_ack;

  reg [15:0] reg_start_address;
  assign start_address = reg_start_address;

  wire frame_receive_error;

  wire frame_received_start_address;
  wire [15:0] frame_start_address_received;

  wire [15:0] frame_remote_address;
  wire  [7:0] frame_remote_length;

  parameter[3:0]
    RECEIVER_IDLE            = 4'b0000,
    SETUP_NEXT_FRAME_RECEIVE = 4'b0001,
    RECEIVING_FRAME          = 4'b0010,
    CANCEL_FRAME_RECEIVE     = 4'b0011,
    WAITING_FOR_ACK_N        = 4'b0100,
    FINALIZE                 = 4'b0101;

  reg [3:0] reg_receiver_state;
  reg [3:0] reg_receiver_next_state;

  reg reg_received_valid_start_frame;

  //
  // Create receiver instance
  //
  menlo_babelfish_rdma_frame_receiver rdma_frame_receiver (
    .fpga_clock(fpga_clock),
    .gigatron_clock(gigatron_clock),
    .reset(reset),

    .famicom_pulse(famicom_pulse),    // hsync_n, famicom_pulse
    .famicom_latch(famicom_latch),    // vsync_n, famicom_latch
    .famicom_data(famicom_data),      // famicom_data

    .request(reg_receive_frames_request),
    .request_ack(receive_frames_request_ack),

    .frame_remote_address(frame_remote_address),
    .frame_remote_length(frame_remote_length),

    .receiver_state(receiver_realtime_state),

    .receive_error(frame_receive_error),
    .receive_error_state(frame_receiver_error_state), // output [4:0]

    .received_start_address(frame_received_start_address),
    .start_address(frame_start_address_received),

    .ram_address(ram_address),
    .ram_data(ram_data),
    .ram_write(ram_write)
  );

  //
  // The receiver is an IDLE state until the receiver request
  // is asserted.
  //
  // It then goes into a receiving frames state and attempts
  // to receive frames until a valid start address frame is received,
  // or the request is de-asserted.
  //
  // Note that since there is no explicit sync as to when reception
  // of a valid frame sequence is to begin a series of attempted frame receives
  // may return errors due to bad a checksum on the frame, as this is just the
  // input data line not yet containing valid frame data.
  //
  // Since each frame starts its receive on the vsync_n rising edge
  // (famicom_latch), this aligns the bit stream with a valid sequence
  // when it starts. Since this is a one way protocol, future checksum
  // errors can't be communicated to the sender.
  //
  // In this logic, checksum errors are accepted until the first valid
  // frame is received. At this point future checksum errors cause reception
  // to stop and an error returned to the caller since one, or more of
  // the programs RDMA transfers will be missing.
  //

  always@(posedge fpga_clock) begin

    if (reset == 1'b1) begin
      reg_receiver_state <= RECEIVER_IDLE;
      reg_receiver_next_state <= RECEIVER_IDLE;
      reg_request_ack <= 1'b0;

      reg_receive_error <= 1'b0;
      reg_receive_error_state <= 0;
      reg_received_valid_start_frame <= 1'b0;
      reg_receive_frames_request <= 1'b0;
      reg_start_address <= 16'h0000;
    end
    else begin

      //
      // Not reset
      //

      case (reg_receiver_state) 
        RECEIVER_IDLE: begin

            if (request == 1'b1) begin

              // These variables track a series of RDMA frame transfers
              reg_receive_error <= 1'b0;
              reg_receive_error_state <= 0;
              reg_received_valid_start_frame <= 1'b0;
              reg_start_address <= 16'h0000;

              reg_receiver_state <= SETUP_NEXT_FRAME_RECEIVE;
            end
        end

        SETUP_NEXT_FRAME_RECEIVE: begin
          reg_receive_frames_request <= 1'b1;
          reg_receiver_state <= RECEIVING_FRAME;
        end

        CANCEL_FRAME_RECEIVE: begin
          // Cancel a frame receive due to an error
          reg_receive_frames_request <= 1'b0;

          // reg_receiver_next_state is set by invoker

          reg_receiver_state <= WAITING_FOR_ACK_N;
        end

        RECEIVING_FRAME: begin

          if (receive_frames_request_ack == 1'b1) begin

              //
              // RDMA frame receiver has ackknowledged the transfer
              //
	      if (frame_receive_error == 1'b1) begin
    
                //
                // The received frame has indicated an error
                //
    
    		if (reg_received_valid_start_frame == 1'b1) begin

		  //
		  // A frame receive error after a valid start frame
		  // is a receiver error to the caller.
		  //

		  // Capture and post the error
		  reg_receive_error_state <= frame_receiver_error_state;
		  reg_receive_error <= 1'b1;

		  // indicate complete to the invoker
		  reg_request_ack <= 1'b1;

		  // Go to FINALIZE state after frame transfer is cancelled
		  reg_receiver_next_state <= FINALIZE;

		  // Cancel frame transfer
		  reg_receiver_state <= CANCEL_FRAME_RECEIVE;
		end
		else begin

		  //
		  // A receive frame error has occurred, but we have not
		  // started a series of RDMA transfers, so this error will
		  // be ignored. Reset the frame receiver for the next
		  // frame synchronization interval.
		  //
		  reg_receiver_next_state <= RECEIVER_IDLE;
		  reg_receiver_state <= CANCEL_FRAME_RECEIVE;
		end
	      end
	      else begin

		//
		// Received a valid frame without error
		//
		if (reg_received_valid_start_frame == 1'b0) begin

		  //
		  // Received valid frame, no more errors allowed till successful
		  // start address frame is received.
		  //
		  reg_received_valid_start_frame <= 1'b1;
		end

		//
		// See if its a start address frame, which ends a series
		// of transfers.
		//
		if (frame_received_start_address == 1'b1) begin

    		  reg_start_address <= frame_start_address_received;

		  // Cancel frame receive
		  reg_receive_frames_request <= 1'b0;

		  // indicate complete to the invoker
		  reg_request_ack <= 1'b1;

		  // Go to FINALIZE state after frame transfer handshake
		  reg_receiver_next_state <= FINALIZE;

		  reg_receiver_state <= WAITING_FOR_ACK_N;
		end
		else begin

		  //
		  // Setup for the next frame receive
		  //
    
    		  // Cancel current frame receive
		  reg_receive_frames_request <= 1'b0;

    		  reg_receiver_next_state <= SETUP_NEXT_FRAME_RECEIVE;

    		  reg_receiver_state <= WAITING_FOR_ACK_N;

		end // next frame receive

	      end // valid frame received

          end // receive_frames_request_ack

        end // end case RECEIVING_FRAME

        WAITING_FOR_ACK_N: begin
          if (receive_frames_request_ack == 1'b0) begin
            // ack has dropped.

            // loader_next_state was set by state receiving the frame.
            reg_receiver_state <= reg_receiver_next_state;
          end
        end

        FINALIZE: begin
          // Stay in finalize state until request is deasserted.
          if (request == 1'b0) begin
            reg_request_ack <= 1'b0;
            reg_receiver_state <= RECEIVER_IDLE;
          end
        end

        default: begin
          reg_receiver_state <= RECEIVER_IDLE;
        end

      endcase

    end // not reset
  end // always

endmodule

//
// Gigatron frame receiver.
//
// The Gigatron frame receiver can be though of as a form of RDMA
// (Remote Direct Memory Access), as each Gigatron frame is a request to
// write a specific memory address, and length in the Gigatrons
// RAM by the loader.
//
// Each RDMA frame can be a subset of a larger memory transfer, tracked by
// the higher level loader based on its loader protocol.
//
// The Gigatron loader frame consists of up to 518 bits which starts sending
// during the end of the VSYNC interval, and clocks each bit at the end of
// the HSYNC interval. This way the bits are sent during the blanking times
// of a VGA monitor.
//
// The frame contains the remote Gigatron memory load address for the data
// portion of the frame, a 6 bit length, and up to 60 bytes of data and a
// checksum.
//
// Frame addresses and length do not cross Gigatron page (256 bytes) boundaries.
//
// A scatter/gather list of loader memory addresses is represented as multiple
// frames sent in sequence, with a last one wins model in regards to any
// memory overlaps.
//
// A received frame length of 0 indicates that its a start program address frame.
//
// If this type of frame is received, its indicated in the output signals, and it
// has no data payload.
//
// The data portion of the received frame is stored in the RAM starting at the
// received remote Gigatron memory address specified in the frame.
//
// The frame's received remote address and length are passed in the output
// signals to the invoker after the data transfer is done.
//
// Frame receive errors are indicated in the error output signals, including
// the state machines value for diagnostics.
//
module menlo_babelfish_rdma_frame_receiver
(
    input fpga_clock,      // FPGA 50Mhz clock
    input gigatron_clock,  // 6.25 Mhz Gigatron clock
    input reset,           // Reset when == 1

    // pulse and latch are the input timing control signals.
    input  famicom_pulse,
    input  famicom_latch,

    // Serial data input
    input  famicom_data,

    // Parameters from BabelFish page receiver state machine.
    input  request,     // frame send request
    output request_ack, // frame send done.

    //
    // This address and length are the values received from the loader frame
    // and represent the remote page address and length.
    //
    output [15:0] frame_remote_address,
    output [7:0]  frame_remote_length,

    //
    // This is a real time indication of the receiver state.
    //
    // bits [3:0] frame state.
    // bits [7:5] bit serializer state.
    //
    output [7:0]  receiver_state,

    // Receive error, and diagnostic state
    output        receive_error,
    output [4:0]  receive_error_state,

    // This indicates if a start address frame is recieved
    output        received_start_address,
    output [15:0] start_address,

    // These are the signals to write bytes to the RAM
    output [15:0] ram_address,
    output [7:0]  ram_data,
    output        ram_write
);

  reg reg_request_ack;
  assign request_ack = reg_request_ack;

  reg reg_received_start_address;
  assign received_start_address = reg_received_start_address;

  reg [15:0] reg_start_address;
  assign start_address = reg_start_address;

  reg [15:0] reg_frame_remote_address;
  assign frame_remote_address = reg_frame_remote_address;

  reg [7:0] reg_frame_remote_length;
  assign frame_remote_length = reg_frame_remote_length;

  reg reg_receive_error;
  assign receive_error = reg_receive_error;

  reg [4:0] reg_receive_error_state;
  assign receive_error_state = reg_receive_error_state;

  // This allows real time monitoring of the bit receiver
  wire [2:0] bit_receiver_state;

  // Loader state machine
  reg [4:0] loader_state;
  reg [4:0] loader_next_state;

  assign receiver_state [4:0] = loader_state;
  assign receiver_state [7:5] = bit_receiver_state;

  reg [15:0] reg_ram_address;
  assign ram_address = reg_ram_address;

  reg [7:0] reg_ram_data;
  assign ram_data = reg_ram_data;

  reg       reg_ram_write;
  assign ram_write = reg_ram_write;

  // Running checksum of the current frame
  reg [7:0] loader_checksum;

  reg [7:0] reg_running_checksum;
  reg [7:0] reg_running_checksum_page;

  //
  // Each frame may be the start of a new page, but we don't
  // know until we get the high address byte. So a running checksum
  // candidate is kept up to date until we receive the high address
  // byte. If the page address has changed, it becomes the new
  // running checksum.
  //
  // In addition, sometimes two back to back GT1 pages contain
  // the same page address, but the loader still resets the checksum
  // for each page. Since we don't have insight into the loaders
  // state the running_checksum_candidate is kept up to date
  // with the start frame as if new page has started. If the final
  // checksum does not compare, the checksum_candidate is compared,
  // and if its correct for the frame checksum, then it becomes
  // the new running checksum for further frames. This models
  // the undisclosed (by the protocol) internal state of the
  // transmitter.
  //
  // Note: The protocol is not modified since its intention is
  // to work with the loader protocol contained inside the binary
  // ROM image for the Gigatron.
  //
  reg [7:0] reg_running_checksum_candidate;

  // Used for shifted frame start byte
  reg [7:0] shifted_frame_start;

  //
  // This indicates when bits are to be sent, the parameters, and the ack.
  //
  reg       reg_receive_bits_request;
  reg       reg_receive_bits_frame_start;
  reg [3:0] reg_receive_bits_count;

  wire [7:0] receive_bits_value;
  wire       receive_bits_request_ack;

  //
  // Receiver States:
  //

  // rdma_frame_receiver states
  parameter[4:0]
    RECEIVE_IDLE            = 5'b00000,
    RECEIVING_START         = 5'b00001, // (command byte) // 8 bits 'L'
    RECEIVING_LENGTH        = 5'b00010, // 6 bits
    RECEIVING_ADDRESS_HIGH  = 5'b00011, // 8 bits
    RECEIVING_ADDRESS_LOW   = 5'b00100, // 8 bits
    RECEIVING_DATA          = 5'b00101, // rom_length 8 bit data bytes
    RECEIVING_CHECKSUM      = 5'b00110, // 8 bits
    RECEIVING_BYTE          = 5'b00111,
    WAITING_FOR_ACK_N       = 5'b01000,
    WRITE_BYTE_TO_RAM       = 5'b01001,
    WRITING_BYTE_TO_RAM     = 5'b01010,
    BYTE_WRITTEN_TO_RAM     = 5'b01011,
    FINALIZE                = 5'b01100,
    SETUP_RAM_TRANSFER      = 5'b01101,
    RECEIVE_NEXT_DATA_BYTE  = 5'b01110,
    RECEIVE_DATA_COMPLETE   = 5'b01111,
    ADDING_SHIFTED_START    = 5'b10000,
    LAST_UNUSED             = 5'b10001;

  // Count of data to receive
  reg [7:0] reg_data_to_receive;

  // total frames received. Wraps around. For debugging/tracing.
  reg [15:0] reg_total_frames_received;

  // Count of error frames
  reg [15:0] reg_total_frames_received_error;

  // Count of checksum error frames
  reg [15:0] reg_total_frames_received_checksum_error;

  //
  // This RDMA implementation uses the BabelFish loaders link layer
  // protocol which is a serial based link layer, with explicit
  // frame timing signals.
  //
  menlo_babelfish_rdma_linklayer_byte_receiver rdma_byte_receiver (
    .fpga_clock(fpga_clock),
    .reset(reset),
    .value(receive_bits_value),
    .number_of_bits(reg_receive_bits_count),
    .pulse(famicom_pulse),          // hsync_n, famicom_pulse
    .latch(famicom_latch),          // vsync_n, famicom_latch
    .frame_start(reg_receive_bits_frame_start),    // set if this is the first byte of the frame.
    .input_port(famicom_data),     // famicom_data
    .receiver_state(bit_receiver_state),
    .request(reg_receive_bits_request),
    .request_ack(receive_bits_request_ack)
  );

  //
  // debug signals
  //
  reg debug_receiving_checksum;

  always@(posedge fpga_clock) begin

    if (reset == 1'b1) begin
      reg_request_ack <= 0;

      reg_frame_remote_address <= 0;
      reg_frame_remote_length <= 0;

      reg_receive_error <= 0;
      reg_receive_error_state <= RECEIVE_IDLE; // 0

      reg_ram_address <= 0;
      reg_ram_data <= 0;
      reg_ram_write <= 0;

      loader_state <= RECEIVE_IDLE;
      loader_next_state <= RECEIVE_IDLE;

      reg_running_checksum <= 0;
      reg_running_checksum_candidate <= 8'h67; // 'g'
      reg_running_checksum_page <= 8'hFF;

      loader_checksum <= 0;

      reg_data_to_receive <= 0;

      shifted_frame_start <= 0;

      reg_received_start_address <= 1'b0;
      reg_start_address <= 0;

      reg_total_frames_received <= 0;
      reg_total_frames_received_error <= 0;
      reg_total_frames_received_checksum_error <= 0;

      //
      // communication variable with the receive bits process.
      //
      reg_receive_bits_request <= 1'b0;
      reg_receive_bits_frame_start <= 1'b0;
      reg_receive_bits_count <= 4'b0;

      //
      // Debug
      //
      debug_receiving_checksum <= 0;

    end
    else begin

      //
      // Not reset
      //

      case (loader_state) 

        RECEIVE_IDLE: begin

          debug_receiving_checksum <= 1'b0;

          if (request == 1'b1) begin

            //
            // Request to receive a frame.
            //
            reg_request_ack <= 0;

            reg_receive_error <= 1'b0;

            reg_total_frames_received <= reg_total_frames_received + 1;

            //
            // checksum starts with 'g' 0x67.
            //
            loader_checksum <= 8'h67;

            reg_running_checksum_candidate <= 8'h67; // 'g'

            shifted_frame_start <= 0;

            // Start byte is 8 bits
            reg_receive_bits_count <= 4'd8;

            //
            // This is the start of a frame.
            //
            // The byte receiver will wait for:
            //
            // vsync_n == HIGH
            //
            // transmitter drives the first bit onto the famicom_data port
            //
            // vsync_n == LOW (negative edge)
            //
            // enters the per bit state machine with hsync_n LOW => HIGH
            // to sample bit.
            //
            reg_receive_bits_frame_start <= 1'b1;

            // Request the bit receiver to go
            reg_receive_bits_request <= 1'b1;

            // return to RECEIVING_START state when done
            loader_next_state <= RECEIVING_START;

            // In RECEIVING_BYTE state
            loader_state <= RECEIVING_BYTE;
          end // request == 1'b1

        end // RECEIVER_IDLE

        RECEIVING_START: begin

          //
          // receive start byte has completed, this is not set for
          // the rest of the bytes.
          //
          reg_receive_bits_frame_start <= 1'b0;

          // Expect first byte with frame_start attribute
          if (receive_bits_value != 8'h4C) begin

            //
            // not start byte 'L' as expected
            //

            reg_total_frames_received_error <= reg_total_frames_received_error + 1;

            if (receive_bits_value == 8'h00) begin

              //
              // We can get 0's during a frame in which no data is sent.
              //
              // In this case go back to the idle state.
              //

              loader_state <= RECEIVE_IDLE;
            end
            else begin

              // Set error, ack invoker, wait in finalize for request de-assert.
              reg_receive_error <= 1'b1;
              reg_receive_error_state <= loader_state;
              reg_request_ack <= 1'b1;
              loader_state <= FINALIZE;
            end
          end
          else begin

            //
            // Got expected start character 0x4C 'L'
            //

            //
            // Note: protocol characters are not written to the RAM, just
            // data.
            //

            //
            // Length is sent as 6 bits in the frame protocol, so only setup
            // to receive 6 bits for length.
            //
            reg_receive_bits_count <= 4'd6;

            //
            // Keep frame checksum updated with each byte received.
            //
            loader_checksum <= loader_checksum + receive_bits_value;

            reg_running_checksum <= 
              reg_running_checksum + receive_bits_value;

            reg_running_checksum_candidate <= 
              reg_running_checksum_candidate + receive_bits_value;

            //
            // Gigatron BabelFish.ino additionally adds the shifted
            // value of the frame start byte to the checksum again.
            //
            shifted_frame_start <= receive_bits_value << 6;

            // Start receive bits in parallel with checksum add.
            reg_receive_bits_request <= 1'b1;

            loader_state <= ADDING_SHIFTED_START;
            end

        end

        ADDING_SHIFTED_START: begin

          // shifted frame start calculation is now available.
          loader_checksum <= loader_checksum + shifted_frame_start;

          reg_running_checksum <= reg_running_checksum + shifted_frame_start;

          reg_running_checksum_candidate <= 
            reg_running_checksum_candidate + shifted_frame_start;

          // Enter receive state
          loader_next_state <= RECEIVING_LENGTH;
          loader_state <= RECEIVING_BYTE;
        end

        RECEIVING_LENGTH: begin

          reg_frame_remote_length <= receive_bits_value;

          // Add the received length byte to the checksum.
          loader_checksum <= loader_checksum + receive_bits_value;

          reg_running_checksum <= 
            reg_running_checksum + receive_bits_value;

          reg_running_checksum_candidate <= 
            reg_running_checksum_candidate + receive_bits_value;

          // The rest of the byte transfers in the frame will be 8 bit.
          reg_receive_bits_count <= 4'd8;

          reg_receive_bits_request <= 1'b1;

          loader_next_state <= RECEIVING_ADDRESS_HIGH;
          loader_state <= RECEIVING_BYTE;
        end

        RECEIVING_ADDRESS_HIGH: begin

          // receive the high address byte
          reg_frame_remote_address[15:8] <= receive_bits_value;

          //
          // If reg_frame_remote_address[15:8] is different
          // than the one we have for the current running checksum
          // it gets reset to its initial value as this
          // represents a new page.
          //
          if (receive_bits_value != reg_running_checksum_page) begin

              reg_running_checksum_page <= receive_bits_value;

              //
              // The running checksum is updated with the candidate.
              //
              reg_running_checksum <= 
                reg_running_checksum_candidate + receive_bits_value;

          end
          else begin

            //
            // Still within the same page, so keep current running checksum
            //
            reg_running_checksum <= 
              reg_running_checksum + receive_bits_value;
          end

          reg_running_checksum_candidate <= 
            reg_running_checksum_candidate + receive_bits_value;

          loader_checksum <= loader_checksum + receive_bits_value;

          reg_receive_bits_request <= 1'b1;

          loader_next_state <= RECEIVING_ADDRESS_LOW;
          loader_state <= RECEIVING_BYTE;
        end

        RECEIVING_ADDRESS_LOW: begin

          // Received the low address byte
          reg_frame_remote_address[7:0] <= receive_bits_value;

          loader_checksum <= loader_checksum + receive_bits_value;

          reg_running_checksum <= reg_running_checksum + receive_bits_value;

          reg_running_checksum_candidate <= 
            reg_running_checksum_candidate + receive_bits_value;

          //
          // reg_frame_remote_length is the total data length
          // to transfer for the current frame.
          //
          // If a length of 0 is received, its a start address frame
          // with zero length data. The start address after reception
          // is returned separately in an output variable/signal to
          // the invoker as its not written to the RAM.
          //
          if (reg_frame_remote_length == 8'h00) begin

              //
              // Start frame. There are no data bytes to receive.
              // Receive the checksum, validate, and set the
              // start address output signal, and complete.
              //
              reg_data_to_receive <= 8'h00;

              // Indicate we received the start address frame
              reg_start_address <= reg_frame_remote_address;
              reg_received_start_address <= 1'b1;

              // Checksum state will set output error if invalid.
              debug_receiving_checksum <= 1'b1;

              reg_receive_bits_request <= 1'b1;

              loader_next_state <= RECEIVING_CHECKSUM;
              loader_state <= RECEIVING_BYTE;
          end
          else begin

              //
              // Begin receiving data bytes and placing into the RAM.
              //

              // Initialize bytes to receive count down
              reg_data_to_receive <= reg_frame_remote_length;

              loader_state <= SETUP_RAM_TRANSFER;
          end
        end

        SETUP_RAM_TRANSFER: begin

          //
          // This is the startup of the RAM transfer for byte 0.
          //

          // Set ram base address from frames remote (memory) address
          reg_ram_address <= reg_frame_remote_address;

          reg_receive_bits_request <= 1'b1;

          loader_next_state <= RECEIVING_DATA;
          loader_state <= RECEIVING_BYTE;
        end

        RECEIVING_DATA: begin

          //
          // Data byte has been received from the link layer.
          //
          // Update the checksum and write it to RAM.
          //
          reg_ram_data <= receive_bits_value;

          loader_checksum <= loader_checksum + receive_bits_value;

          reg_running_checksum <= reg_running_checksum + receive_bits_value;

          reg_running_checksum_candidate <= 
            reg_running_checksum_candidate + receive_bits_value;

          // Decrement the transfer count to account for the byte.
          reg_data_to_receive <= reg_data_to_receive - 1;

          loader_next_state <= RECEIVE_NEXT_DATA_BYTE;

          // Write the byte to the RAM
          loader_state <= WRITE_BYTE_TO_RAM;
        end

        RECEIVE_NEXT_DATA_BYTE: begin

          //
          // This is for a continuing transfer other than byte 0
          // after the just received byte has been written to RAM.
          //
          if (reg_data_to_receive == 8'h00) begin

            // Checksum state will set output error if invalid.
            debug_receiving_checksum <= 1'b1;

            // Done with data transfer, receive the checksum from the transmitter.
            reg_receive_bits_request <= 1'b1;

            loader_next_state <= RECEIVING_CHECKSUM;
            loader_state <= RECEIVING_BYTE;
          end
          else begin

            // The reg_data_to_receive count has already been decremented

            // Advance the RAM address
            reg_ram_address <= reg_ram_address + 1;

            reg_receive_bits_request <= 1'b1;

            loader_next_state <= RECEIVING_DATA;
            loader_state <= RECEIVING_BYTE;
          end
        end

        RECEIVING_CHECKSUM: begin

          //
          // Validate the check sum is what is expected.
          //
          // TODO: validating...
          //if (receive_bits_value != loader_checksum) begin

          if ((receive_bits_value + reg_running_checksum) != 8'h00) begin

            //
            // This may be a start of a new page with the same
            // page address as a previous one.
            //
            if ((receive_bits_value + reg_running_checksum_candidate) != 8'h00) begin

              // Set error, ack invoker, wait in finalize for request de-assert.
              reg_receive_error <= 1'b1;
              reg_receive_error_state <= loader_state;

              reg_total_frames_received_error <= reg_total_frames_received_error + 1;

              reg_total_frames_received_checksum_error <= 
                reg_total_frames_received_checksum_error + 1;
            end
            else begin

              //
              // Make the current running checksum the candidate so future
              // frames will be received correctly.
              //
              reg_running_checksum <= reg_running_checksum_candidate;
            end
          end

          loader_state <= RECEIVE_DATA_COMPLETE;
        end

        RECEIVE_DATA_COMPLETE: begin

          // Done with frame, checksum is valid
          reg_request_ack <= 1'b1;

          // Finalize waits for request to deassert
          loader_state <= FINALIZE;
        end

        FINALIZE: begin

          // Stay in finalize state until request is deasserted.
          if (request == 1'b0) begin
            reg_request_ack <= 1'b0;
            loader_state <= RECEIVE_IDLE;
          end

        end

        //
        // Reading a byte from the ROM and then sending it to the
        // babelfish_bit_sender is a common operation used for
        // each byte in the frame envelope, so make it a common
        // state machine.
        //

        WRITE_BYTE_TO_RAM: begin

          //
          // reg_ram_address, reg_ram_data, loader_next_state
          // has been set by invoker.
          //
          // This entry gives 1 clock to access RAM
          //

          reg_ram_write <= 1'b1;

          loader_state <= WRITING_BYTE_TO_RAM;
        end

        WRITING_BYTE_TO_RAM: begin
          // byte in reg_ram_data stored in ram

          reg_ram_write <= 1'b0;

          // 1 clock delay for deassert of reg_ram_write
          loader_state <= BYTE_WRITTEN_TO_RAM;
        end

        BYTE_WRITTEN_TO_RAM: begin
          loader_state <= loader_next_state;
        end

        //
        // Each byte received uses the following two states to handle
        // hand shake with the babelfish_bit_receiver module.
        //
        // loader_next_state is used to return to the previous transfer
        // phase when done.
        //

        RECEIVING_BYTE: begin
          // Receiving byte. Wait for ACK from byte receiver.
          if (receive_bits_request_ack == 1'b1) begin
            // Request has acknowledged, deassert request, wait for ack to drop.
            reg_receive_bits_request <= 1'b0;
            loader_state <= WAITING_FOR_ACK_N;
          end
        end

        WAITING_FOR_ACK_N: begin
          if (receive_bits_request_ack == 1'b0) begin
            // ack has dropped.

            // loader_next_state was set by state receiving the byte.
            loader_state <= loader_next_state;
          end
        end

        default: begin
          loader_state <= RECEIVE_IDLE;
        end

      endcase

    end

  end // always

  //
  // The Gigatron/BabelFish frame protocol is as follows:
  //
  // A bit stream of 518 total bits.
  //
  // Start of the bitstream is clocked by gigatron_famicom_latch (vsync_n) going high.
  //
  // Each bit is clocked by gigatron_famicom_pulse (hsync_n) going high.
  //
  // The bit is placed on gigatron_famicom_data as input to the Gigatron.
  // 
  // Order sent:
  //
  // Note: all bits are sent MSB first.
  //
  // 8 bits - start byte 'L' (0x4C)
  // 6 bits - block_length
  // 8 bits - address_high
  // 8 bits - address_low
  // 8 bits - data_byte[0]
  // 8 bits - data_byte [block_length - 1]
  // 8 bits - checksum
  //
  
  //
  // Note: There is a place where (2) bits are dropped on purpose
  // due to Gigatron loader timings. Ensure this is implemented
  // in the state machine above. It shows up in the (6) bit
  // length period.
  //

endmodule // menlo_babelfish_frame_receiver

//
// RDMA Link Layer Byte Receiver for Gigatron BabelFish Protocol.
//
// This implementation uses the Gigatron BabelFish serial loader
// protocol and signals for implementation. Other RDMA LinkLayer
// receivers would have different framing models, such as
// ethernet/ip packets.
//
// Receive bits from the input port.
//
// latch is the vsync_n signal from the Gigatron which indicates
// the start of the frame to receive.
//
// pulse is the hsync_n signal from the Gigatron which times
// the bit send rate from the transmitter.
//
// frame_start is set for the first byte of the frame and syncs
// with vsync_n (latch) before receiving the rest of the frame. It
// should only be set for the first byte of the frame, and only
// the first bit will wait for vsync_n transition.
//
// Bits are sent MSB first, up to number_of_bits.
//
// Since the Gigatron frame protocol uses a variable number
// of bits without an explicit start/stop signal for character
// frames, the number of bits expected are passed by the invoker,
// which implements the RDMA receive frame state machine.
//
// Request handshake protocol:
//
// See menlo_babelfish_bit_sender.
//
// Receiver: (this module implementing the RDMA receiver)
//
// Receiver starts with request and request_ack == 1'b0 and
// internally in the IDLE state.
//
// Receiver when in IDLE state receives request == 1'b1, and sets
// an internal register to latch the request. It then performs the
// request asynchronously based on its internal state machine.
//
// When the request is complete it sets request_ack == 1'b1, and
// then goes into a state to await the de-assertion of request to 1'b0.
//
// When request becomes 1'b0, it clears request_ack and goes back
// to the idle state to begin await a new request.
//
module menlo_babelfish_rdma_linklayer_byte_receiver (
  input fpga_clock,
  input reset,          // high true
  output [7:0] value,   // received value.
  input [3:0] number_of_bits, // number of bits in the byte frame.
  input pulse,          // hsync_n, famicom_pulse
  input latch,          // vsync_n, famicom_latch
  input frame_start,    // set if this is the first byte of the frame.
  input input_port,     // famicom_data
  output [2:0] receiver_state, // exposed receiver state
  input  request,
  output request_ack
  );

  reg [7:0] reg_receive_bits_value;
  assign value = reg_receive_bits_value;

  reg reg_request_ack;
  assign request_ack = reg_request_ack;

  //
  // state is exposed to the caller to allow it to monitor
  // the transfer in case of errors, timeout, etc.
  //
  // A reset clears the receiver for a restart.
  //
  // This module does not impose a timeout, but exposes
  // its state for the invoker to determine.
  //
  reg [2:0] bits_state;
  assign receiver_state = bits_state;

  // rdma_byte_receiver states
  parameter[2:0]
    BITS_IDLE               = 3'b000,
    BITS_TRANSFER_BIT       = 3'b001,
    BITS_WAIT_H_PULSE_LOW   = 3'b010,
    BITS_WAIT_H_PULSE_HIGH  = 3'b011,
    BITS_WAIT_V_LATCH_LOW   = 3'b100,
    BITS_WAIT_V_LATCH_HIGH  = 3'b101,
    BITS_SENDING_ACK        = 3'b110,
    BITS_UNASSIGNED         = 3'b111;

  // Bits are sent MSB first, so this counts down.
  reg [3:0] reg_bits_counter;

  // total bytes received. Wraps around. For debugging/tracing.
  reg [15:0] reg_total_bytes_received;

  always@(posedge fpga_clock) begin

    if (reset == 1'b1) begin
      reg_receive_bits_value <= 0;
      reg_request_ack <= 1'b0;
      bits_state <= BITS_IDLE;
      reg_bits_counter <= 1'b0;
      reg_total_bytes_received <= 0;
    end
    else begin

      //
      // Not reset
      //

      case (bits_state) 

        BITS_IDLE: begin

          if (request == 1'b1) begin

            //
            // Command to receive count bits into the value register.
            //

            //
            // Sequence is bit number 7 - 0 for 8 bit, and 5 - 0 for 6 bit receive.
            //
            reg_bits_counter <= number_of_bits - 1;

            reg_receive_bits_value <= 0;

            reg_total_bytes_received <= reg_total_bytes_received + 1;

            if (frame_start == 1'b1) begin

              //
              // First bit of first byte syncs with vsync_n for start of frame.
              //
              // Frame start sequence:
              //
              // 1) Receiver waits for vsync_n to be HIGH
              //
              // 2) Transmitter drives first bit onto output port
              //
              // 3) Receiver waits for vsync_n going LOW (negative edge)
              //
              // Note: At his point its the normal per bit handshake
              // with hsync_n.
              //
              // 4) Receiver waits for hsync_n to be LOW
              //
              // 5) Receiver waits for hsync_n to be HIGH (positive edge)
              //
              // 6) Receiver samples the data at this edge.
              //
              // 7) Receive rest of 7 bits using normal per bit handshake.
              //
              bits_state <= BITS_WAIT_V_LATCH_HIGH;
            end
            else begin
              bits_state <= BITS_TRANSFER_BIT;
            end

          end
        end

        BITS_TRANSFER_BIT: begin

          //
          // Note end is underflow wrap around since bit 0 must be received.
          //
          if (reg_bits_counter != 4'b1111) begin
            bits_state <= BITS_WAIT_H_PULSE_LOW;
          end
          else begin
            reg_request_ack <= 1'b1;
            bits_state <= BITS_SENDING_ACK;
          end
        end

        BITS_WAIT_H_PULSE_LOW: begin

          //
          // Waiting for pulse to be low
          //
          if (pulse == 1'b0) begin
            bits_state <= BITS_WAIT_H_PULSE_HIGH;
          end
        end

        BITS_WAIT_H_PULSE_HIGH: begin

          //
          // Waiting for pulse to be high
          //
          if (pulse == 1'b1) begin

            //
            // The input port is sampled on the rising edge of hsync_n going HIGH.
            //
            reg_receive_bits_value[reg_bits_counter] <= input_port;
            reg_bits_counter <= reg_bits_counter - 1;

            // Back to transfer next bit
            bits_state <= BITS_TRANSFER_BIT;
          end
        end

        BITS_WAIT_V_LATCH_HIGH: begin

          //
          // Waiting for vsync_n latch signal to be HIGH
          //
          if (latch == 1'b1) begin

            //
            // vsync_n is HIGH, which arms the frame start sequence.
            //
            // Wait for vsync_n LOW before starting the frame receive.
            //

            bits_state <= BITS_WAIT_V_LATCH_LOW;
          end
        end

        BITS_WAIT_V_LATCH_LOW: begin

          //
          // Waiting for sync_n latch signal to be low
          //
          if (latch == 1'b0) begin

            //
            // The frame receive has begin. Enter the bits transfer
            // handshake state.
            //
            bits_state <= BITS_TRANSFER_BIT;
          end
        end

        BITS_SENDING_ACK: begin

          //
          // Waiting for request to be de-asserted
          //
          if (request == 1'b0) begin
            reg_request_ack <= 1'b0;
            bits_state <= BITS_IDLE;
          end

        end

        default: begin
        end

      endcase

    end // not reset

  end // always sendBits

endmodule // menlo_babelfish_bit_receiver

//
// Test benches
//
// The following test benches are great not just for validating
// components but for exploring the design. It allows you to update
// the test bench to exercise a specific component and see its exact
// behavior, before and after any modifications.
//

`define tb_menlo_babelfish_assert(signal, value) \
    if (signal !== value) begin \
	     $display("ASSERTION FAILED in %m: signal != value"); \
		  $stop; \
    end

module tb_menlo_babelfish();

  // Validation loop variables
  integer index;
  integer rom_a;
  integer ram_a;

  reg [7:0] rom_value;
  reg [7:0] ram_value;
  reg [7:0] page_length;
  reg [15:0] full_address;

  reg compare_error;

  // FPGA clock
  reg fpga_clock;

  // VGA clock
  reg vga_clock;

  // Gigatron clock
  reg clock_6_25;

  reg reset;

  // VGA signals
  wire hsync_n;
  wire vsync_n;

  // Serial game controller
  wire famicom_pulse;
  wire famicom_latch;

  // The game control pulse, latch is driven by the VGA signals.
  assign famicom_pulse = hsync_n;
  assign famicom_latch = vsync_n;

  // output from transmitter, input to receiver
  wire  famicom_data;

  // transmitter control signals
  reg reg_transmitter_request;
  wire transmitter_request_ack;

  parameter ROM_ARRAY_SIZE = 32767;

  //  width                      depth
  reg [7:0] reg_option_rom_array [0:ROM_ARRAY_SIZE];

  wire [15:0] rom_address;
  reg [7:0]   reg_rom_data;

  //
  // The RAM is loaded by the receiver and its data is analyzed
  // against the ROM images data pages at the end of the test.
  //
  parameter RAM_ARRAY_SIZE = 32767;

  reg [7:0]   reg_ram_array [0:RAM_ARRAY_SIZE];

  wire [15:0] ram_address;
  wire  [7:0] ram_data;
  wire        ram_write;
  reg [7:0]   reg_ram_read_data;

  //
  // This is a comparison RAM used by the testbench
  // after the RDMA transfer of the GT1 file has completed.
  //
  reg [7:0]   reg_compare_ram_array [0:RAM_ARRAY_SIZE];

  // Test control signals
  reg reg_test_done;
  reg reg_receive_error;
  reg reg_receiver_done;
  reg reg_transmitter_done;

  // Device Under Test instance (Transmitter)
  menlo_babelfish_rdma_transmitter rdma_transmitter (
    .fpga_clock(fpga_clock),
    .gigatron_clock(clock_6_25),
    .reset(reset),

    .famicom_pulse(famicom_pulse),
    .famicom_latch(famicom_latch),
    .famicom_data(famicom_data), // output

    .request(reg_transmitter_request),
    .request_ack(transmitter_request_ack),

    .rom_address(rom_address),
    .rom_data(reg_rom_data)
  );

  //
  // RDMA Receiver signals
  //
  reg reg_receiver_request;
  wire receiver_request_ack;

  wire [15:0] received_start_address;

  wire [7:0]  receiver_state;
  wire        receive_error;
  wire [7:0]  receive_error_state;

  // Device Under Test instance (Receiver)
  menlo_babelfish_rdma_receiver rdma_receiver (
    .fpga_clock(fpga_clock),
    .gigatron_clock(clock_6_25),
    .reset(reset),

    .famicom_pulse(famicom_pulse),
    .famicom_latch(famicom_latch),
    .famicom_data(famicom_data), // input

    .request(reg_receiver_request),
    .request_ack(receiver_request_ack),

    .start_address(received_start_address),

    .receiver_realtime_state(receiver_state),

    .receive_error(receive_error),
    .receive_error_state(receive_error_state),

    .ram_address(ram_address),
    .ram_data(ram_data),
    .ram_write(ram_write)
  );

  //
  // Video sync generator instance
  //
  wire blank_n;

  video_sync_generator video_signal_generator(
    .reset(reset),
    .vga_clk(vga_clock),
    .blank_n(blank_n),
    .HS(hsync_n),
    .VS(vsync_n)
  );

  // Set initial values
  initial begin

     // Validation loop variables
     index = 0;
     rom_a = 0;
     ram_a = 0;
     rom_value = 0;
     ram_value = 0;
     page_length = 0;
     full_address = 0;
     compare_error = 0;

     fpga_clock = 0;
     vga_clock = 0;
     clock_6_25 = 0;
     reset = 1;
     reg_transmitter_request = 0;
     reg_receiver_request = 0;

     // Test control signals
     reg_test_done = 0;
     reg_receive_error = 0;
     reg_receiver_done = 0;
     reg_transmitter_done = 0;

     //
     // tetris.gt1 binary rom image file converted with:
     //
     // hexdump -v  -e '1/1  "%02X\n"' tetris.gt1 >gt1_tetris_verilog_data.txt
     //

     reg_rom_data = 0;

     $readmemh(
       "C:/Dropbox/embedded/altera/workspace/menlo_gigatron_de10_nano/gt1_tetris_verilog_data.txt",
        reg_option_rom_array
       );

    reg_ram_read_data = 0;

    //
    // Initialize the RAM contents
    //
    for (index = 0; index < RAM_ARRAY_SIZE; index = index + 1) begin
      reg_ram_array[index] = 0;
    end

    for (index = 0; index < RAM_ARRAY_SIZE; index = index + 1) begin
      reg_compare_ram_array[index] = 0;
    end

  end

  //
  // Setup FPGA 50Mhz clock
  //
  // 50mhz == 20ns period.
  // #10 delay is 1/2 of the cycle.
  //
  always #10 fpga_clock = ~fpga_clock;

  //
  // Setup 25Mhz VGA clock
  //
  always #20 vga_clock = ~vga_clock;

  //
  // Setup 6.25Mhz Gigatron clock at 1ns resolution in simulation.
  //
  // #xx - delay in nanoseconds
  //
  // 6.25mhz == 160ns per cycle.
  //
  // so #80 delay is 1/2 of the cycle.
  //

  always #80 clock_6_25 = ~clock_6_25;

  //
  // ROM implementation
  //
  always @* begin
    reg_rom_data = reg_option_rom_array[rom_address];
  end

  //
  // RAM implementation
  //
  // ram_data - write data when ram_write == 1'b1
  // reg_ram_read_data - RAM data when ram_write != 1'b1
  //
  // Include ram_address and ram-write in sensitivity list.
  //
  always @* begin
    if (ram_write == 1'b1) begin
      reg_ram_array[ram_address] = ram_data; // output from RDMA receiver
    end
    else begin
      // read side
      reg_ram_read_data = reg_ram_array[ram_address];
    end
  end

  //
  // This process monitors the transfers until completed,
  // or an error indication.
  //

  always @(posedge fpga_clock) begin

    if (reset == 1'b1) begin
      reg_test_done <= 1'b0;
      reg_receive_error <= 1'b0;
      reg_transmitter_done <= 1'b0;
      reg_receiver_done <= 1'b0;
    end
    else begin

        // Indication that the receiver is active
    	if (reg_receiver_request == 1'b1) begin
	  if (receive_error == 1'b1) begin
    	    reg_receive_error <= 1'b1;
            // Receiver is done on error signal
            //reg_receiver_request <= 1'b0;
            reg_receiver_done <= 1'b1;
          end
    
          if (receiver_request_ack == 1'b1) begin
           // Receiver has completed.
    	   reg_receiver_done <= 1'b1;
          end
	end

        // Indication that the transmitter is active
	if (reg_transmitter_request == 1'b1) begin
	  if (transmitter_request_ack == 1'b1) begin
            // Transmitter has completed.
	    reg_transmitter_done <= 1'b1;
	  end
	end

        //
	// Test done when a receive error occurs, or when both the
        // transmitter and receiver complete.
        //
	if ((reg_receive_error) || (reg_transmitter_done && reg_receiver_done)) begin
	  reg_test_done <= 1'b1;
	end

    end // not reset

  end

  // Stimulus to step through values
  initial begin

    // Set Reset
    reset = 1'b1;

    // Wait some Gigatron clock cycles
    @(posedge clock_6_25);
    @(posedge clock_6_25);
    @(posedge clock_6_25);
    @(posedge clock_6_25);

    //
    // The RDMA transmitter sends the contents of the memory
    // pages in the ROM which are described in GT1 file format.
    //
    // The RDMA receiver receives these pages as RDMA frames
    // and writes to the RAM memory at the address, length of
    // each frame.
    //
    // At the end of the test, the GT1 file data in the ROM is
    // compared what is in the RAM.
    //
    // Note: Pages in the GT1 file may overlap, with a last sent
    // wins rule. This must be handled in the test.
    //

    // Remove reset
    reset = 1'b0;

    // Wait some clock cycles
    @(posedge fpga_clock);
    @(posedge fpga_clock);
     
    //
    // Initialize the compare ram array.
    //
    // Sections in GT1 files can overlap, and be seen
    // again. This is allowed with a "last one wins" rule.
    //
    // So an additional compare ram memory is initialized with
    // the GT1 file contents, and then used for the final
    // compare.
    //

    rom_a = 0;
    ram_a = 0;

    for (rom_a = 0; rom_a < ROM_ARRAY_SIZE; rom_a = rom_a + 0) begin

      // Get the high address byte of page record.
      full_address[15:8] = reg_option_rom_array[rom_a];

      // High address byte 0, and not ROM location 0 means end of page records.
      if ((full_address[15:8] == 8'h00) && (rom_a != 0)) begin
        // We are done if high_address == 0 not at start of ROM.

        // The start address frame is just after the current 0.
        // Skip 0
        rom_a = rom_a + 1;

        // High start address
        full_address[15:8] = reg_option_rom_array[rom_a];

        rom_a = rom_a + 1;

        // low start address
        full_address[7:0] = reg_option_rom_array[rom_a];
        rom_a = rom_a + 1;

        $display("*** start_address %h", full_address);

        // exit for() loop
        break;
      end

      // Advance past address high byte
      rom_a = rom_a + 1;

      // Address low byte of page
      full_address[7:0] = reg_option_rom_array[rom_a];
      rom_a = rom_a + 1;

      // page length byte
      page_length = reg_option_rom_array[rom_a];
      rom_a = rom_a + 1;

      $display("page remote address %h, length %h", full_address, page_length);

      //
      // Data area in ROM is just after the header above and
      // rom_a points to it.
      //

      // Data area in RAM is the pages specified address
      ram_a = full_address;

      for (index = 0; index < page_length; index = index + 1) begin

        // Get data bytes from the ROM and copy to the RAM.
        rom_value = reg_option_rom_array[rom_a + index];

        reg_compare_ram_array[ram_a + index] = rom_value;

      end // end for data range validate

      // Advance the page data area to the next header start.
      rom_a = rom_a + page_length;

    end // for process GT1 file sections for the compare_ram_array

    // Wait some clock cycles
    @(posedge fpga_clock);
    @(posedge fpga_clock);

    // Set request for receiver first
    reg_receiver_request = 1'b1;

    // Wait some clock cycles
    @(posedge fpga_clock);
    @(posedge fpga_clock);
    @(posedge fpga_clock);
    @(posedge fpga_clock);

    // Set request for transmitter
    reg_transmitter_request = 1'b1;

    @(posedge fpga_clock);
    @(posedge fpga_clock);

    //
    // Wait till test done, or error
    //

    @(posedge reg_test_done);

    // Check for error, stop if so to debug in ModelSim
    if (reg_receive_error == 1'b1) begin
      // Wait two clocks before ending
      @(posedge fpga_clock);
      @(posedge fpga_clock);
      $display("*** RECEIVE ERROR *** Stopped due to reg_receive_error == 1");
      $stop;
    end

    //
    // Note: both transmitter and receiver should be idle here
    // if no error was indicated.
    //

    // Stop transmitter
    reg_transmitter_request = 1'b0;
    @(posedge fpga_clock);
    @(posedge fpga_clock);

    // Stop receiver
    reg_receiver_request = 1'b0;
    @(posedge fpga_clock);
    @(posedge fpga_clock);

    //
    // Compare the output RAM from the receiver with the compare
    // RAM initialized earlier.
    //

    rom_a = 0;
    ram_a = 0;

    for (rom_a = 0; rom_a < ROM_ARRAY_SIZE; rom_a = rom_a + 0) begin

      // Get the high address byte of page record.
      full_address[15:8] = reg_option_rom_array[rom_a];

      // High address byte 0, and not ROM location 0 means end of page records.
      if ((full_address[15:8] == 8'h00) && (rom_a != 0)) begin
        // We are done if high_address == 0 not at start of ROM.

        if (compare_error != 1'b0) begin
            $display("*** FAILED *** RAM contents did not compare to ROM contents for RDMA transfer");
        end
        else begin
            $display("*** PASSED *** RAM contents compare to ROM contents for RDMA transfer");
        end

        // The start address frame is just after the current 0.
        // Skip 0
        rom_a = rom_a + 1;

        // High start address
        full_address[15:8] = reg_option_rom_array[rom_a];

        rom_a = rom_a + 1;

        // low start address
        full_address[7:0] = reg_option_rom_array[rom_a];
        rom_a = rom_a + 1;

        $display("*** start_address %h", full_address);

        $stop;
      end

      // Advance past address high byte
      rom_a = rom_a + 1;

      // Address low byte of page
      full_address[7:0] = reg_option_rom_array[rom_a];
      rom_a = rom_a + 1;

      // page length byte
      page_length = reg_option_rom_array[rom_a];
      rom_a = rom_a + 1;

      $display("page remote address %h, length %h", full_address, page_length);

      //
      // Data area in ROM is just after the header above and
      // rom_a points to it.
      //

      // Data area in RAM is the pages specified address
      ram_a = full_address;

      for (index = 0; index < page_length; index = index + 1) begin

        // Get data bytes from the ROM and compare to the RAM.
        rom_value = reg_option_rom_array[rom_a + index];

        ram_value = reg_ram_array[ram_a + index];

        if (ram_value != rom_value) begin

          $display("*** FAILED *** RAM contents don't match");
          $display("ram_address %h, data %h", ram_a + index, ram_value);
          $display("rom_address %h, data %h", rom_a + index, rom_value);
          $display("May be due to later write, check page addresses of following writes.");

          compare_error <= 1'b1;

          // Let's look at all the pages instead of stopping.
          break;

        end

      end // end for data range validate

      // Advance the page data area to the next header start.
      rom_a = rom_a + page_length;

    end // for process GT1 file sections

    // Wait two clocks before ending
    @(posedge fpga_clock);
    @(posedge fpga_clock);

    $display("*** ERROR *** Ran off end of ROM without termination");

    $stop;

  end // initial

endmodule
